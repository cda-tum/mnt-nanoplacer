module top (
    \A0 , \A1 , \A2 , \A3 , \A4 , \A5 , \A6 , \A7 , \A8 ,
    \A9 , \A10 , \A11 , \A12 , \A13 , \A14 , \A15 , \A16 ,
    \A17 , \A18 , \A19 , \A20 , \A21 , \A22 , \A23 , \A24 ,
    \A25 , \A26 , \A27 , \A28 , \A29 , \A30 , \A31 , \A32 ,
    \A33 , \A34 , \A35 , \A36 , \A37 , \A38 , \A39 , \A40 ,
    \A41 , \A42 , \A43 , \A44 , \A45 , \A46 , \A47 , \A48 ,
    \A49 , \A50 , \A51 , \A52 , \A53 , \A54 , \A55 , \A56 ,
    \A57 , \A58 , \A59 , \A60 , \A61 , \A62 , \A63 , \A64 ,
    \A65 , \A66 , \A67 , \A68 , \A69 , \A70 , \A71 , \A72 ,
    \A73 , \A74 , \A75 , \A76 , \A77 , \A78 , \A79 , \A80 ,
    \A81 , \A82 , \A83 , \A84 , \A85 , \A86 , \A87 , \A88 ,
    \A89 , \A90 , \A91 , \A92 , \A93 , \A94 , \A95 , \A96 ,
    \A97 , \A98 , \A99 , \A100 , \A101 , \A102 , \A103 ,
    \A104 , \A105 , \A106 , \A107 , \A108 , \A109 , \A110 ,
    \A111 , \A112 , \A113 , \A114 , \A115 , \A116 , \A117 ,
    \A118 , \A119 , \A120 , \A121 , \A122 , \A123 , \A124 ,
    \A125 , \A126 , \A127 ,
    \P0 , \P1 , \P2 , \P3 , \P4 , \P5 , \P6 , F  );
  input  \A0 , \A1 , \A2 , \A3 , \A4 , \A5 , \A6 , \A7 ,
    \A8 , \A9 , \A10 , \A11 , \A12 , \A13 , \A14 , \A15 ,
    \A16 , \A17 , \A18 , \A19 , \A20 , \A21 , \A22 , \A23 ,
    \A24 , \A25 , \A26 , \A27 , \A28 , \A29 , \A30 , \A31 ,
    \A32 , \A33 , \A34 , \A35 , \A36 , \A37 , \A38 , \A39 ,
    \A40 , \A41 , \A42 , \A43 , \A44 , \A45 , \A46 , \A47 ,
    \A48 , \A49 , \A50 , \A51 , \A52 , \A53 , \A54 , \A55 ,
    \A56 , \A57 , \A58 , \A59 , \A60 , \A61 , \A62 , \A63 ,
    \A64 , \A65 , \A66 , \A67 , \A68 , \A69 , \A70 , \A71 ,
    \A72 , \A73 , \A74 , \A75 , \A76 , \A77 , \A78 , \A79 ,
    \A80 , \A81 , \A82 , \A83 , \A84 , \A85 , \A86 , \A87 ,
    \A88 , \A89 , \A90 , \A91 , \A92 , \A93 , \A94 , \A95 ,
    \A96 , \A97 , \A98 , \A99 , \A100 , \A101 , \A102 ,
    \A103 , \A104 , \A105 , \A106 , \A107 , \A108 , \A109 ,
    \A110 , \A111 , \A112 , \A113 , \A114 , \A115 , \A116 ,
    \A117 , \A118 , \A119 , \A120 , \A121 , \A122 , \A123 ,
    \A124 , \A125 , \A126 , \A127 ;
  output \P0 , \P1 , \P2 , \P3 , \P4 , \P5 , \P6 , F;
  wire n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147,
    n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159,
    n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
    n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183,
    n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195,
    n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207,
    n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219,
    n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
    n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
    n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255,
    n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267,
    n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
    n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291,
    n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
    n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
    n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327,
    n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339,
    n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351,
    n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
    n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
    n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
    n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
    n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
    n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
    n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
    n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
    n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
    n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
    n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
    n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
    n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
    n508, n509, n510, n512, n513, n514, n515, n516, n517, n518, n519, n520,
    n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
    n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
    n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
    n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
    n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
    n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
    n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
    n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
    n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
    n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
    n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
    n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
    n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
    n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
    n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
    n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
    n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
    n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
    n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
    n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n760, n761,
    n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
    n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
    n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797,
    n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809,
    n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821,
    n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
    n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845,
    n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857,
    n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869,
    n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
    n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
    n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
    n906, n907, n908, n910, n911, n912, n913, n914, n915, n916, n917, n918,
    n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930,
    n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942,
    n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954,
    n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966,
    n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978,
    n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990,
    n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001,
    n1002, n1003, n1004, n1005, n1006, n1007, n1009, n1010, n1011, n1012,
    n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
    n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
    n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
    n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
    n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
    n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
    n1073, n1074, n1075, n1076, n1078, n1079, n1080, n1081, n1082, n1083,
    n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
    n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
    n1104, n1107, n1108, n1109, n1110, n1111, n1112, n1113;
  assign n137 = ~\A125  & \A127 ;
  assign n138 = \A126  & \A127 ;
  assign n139 = \A126  & ~n138;
  assign n140 = \A125  & ~n139;
  assign n141 = ~n137 & ~n140;
  assign n142 = ~\A123  & ~n141;
  assign n143 = ~\A124  & ~n139;
  assign n144 = \A124  & ~n141;
  assign n145 = ~n143 & ~n144;
  assign n146 = \A123  & ~n145;
  assign n147 = ~n142 & ~n146;
  assign n148 = ~\A121  & ~n147;
  assign n149 = ~\A122  & ~n145;
  assign n150 = \A122  & ~n147;
  assign n151 = ~n149 & ~n150;
  assign n152 = \A121  & ~n151;
  assign n153 = ~n148 & ~n152;
  assign n154 = ~\A119  & ~n153;
  assign n155 = ~\A120  & ~n151;
  assign n156 = \A120  & ~n153;
  assign n157 = ~n155 & ~n156;
  assign n158 = \A119  & ~n157;
  assign n159 = ~n154 & ~n158;
  assign n160 = ~\A117  & ~n159;
  assign n161 = ~\A118  & ~n157;
  assign n162 = \A118  & ~n159;
  assign n163 = ~n161 & ~n162;
  assign n164 = \A117  & ~n163;
  assign n165 = ~n160 & ~n164;
  assign n166 = ~\A115  & ~n165;
  assign n167 = ~\A116  & ~n163;
  assign n168 = \A116  & ~n165;
  assign n169 = ~n167 & ~n168;
  assign n170 = \A115  & ~n169;
  assign n171 = ~n166 & ~n170;
  assign n172 = ~\A113  & ~n171;
  assign n173 = ~\A114  & ~n169;
  assign n174 = \A114  & ~n171;
  assign n175 = ~n173 & ~n174;
  assign n176 = \A113  & ~n175;
  assign n177 = ~n172 & ~n176;
  assign n178 = ~\A111  & ~n177;
  assign n179 = ~\A112  & ~n175;
  assign n180 = \A112  & ~n177;
  assign n181 = ~n179 & ~n180;
  assign n182 = \A111  & ~n181;
  assign n183 = ~n178 & ~n182;
  assign n184 = ~\A109  & ~n183;
  assign n185 = ~\A110  & ~n181;
  assign n186 = \A110  & ~n183;
  assign n187 = ~n185 & ~n186;
  assign n188 = \A109  & ~n187;
  assign n189 = ~n184 & ~n188;
  assign n190 = ~\A107  & ~n189;
  assign n191 = ~\A108  & ~n187;
  assign n192 = \A108  & ~n189;
  assign n193 = ~n191 & ~n192;
  assign n194 = \A107  & ~n193;
  assign n195 = ~n190 & ~n194;
  assign n196 = ~\A105  & ~n195;
  assign n197 = ~\A106  & ~n193;
  assign n198 = \A106  & ~n195;
  assign n199 = ~n197 & ~n198;
  assign n200 = \A105  & ~n199;
  assign n201 = ~n196 & ~n200;
  assign n202 = ~\A103  & ~n201;
  assign n203 = ~\A104  & ~n199;
  assign n204 = \A104  & ~n201;
  assign n205 = ~n203 & ~n204;
  assign n206 = \A103  & ~n205;
  assign n207 = ~n202 & ~n206;
  assign n208 = ~\A101  & ~n207;
  assign n209 = ~\A102  & ~n205;
  assign n210 = \A102  & ~n207;
  assign n211 = ~n209 & ~n210;
  assign n212 = \A101  & ~n211;
  assign n213 = ~n208 & ~n212;
  assign n214 = ~\A99  & ~n213;
  assign n215 = ~\A100  & ~n211;
  assign n216 = \A100  & ~n213;
  assign n217 = ~n215 & ~n216;
  assign n218 = \A99  & ~n217;
  assign n219 = ~n214 & ~n218;
  assign n220 = ~\A97  & ~n219;
  assign n221 = ~\A98  & ~n217;
  assign n222 = \A98  & ~n219;
  assign n223 = ~n221 & ~n222;
  assign n224 = \A97  & ~n223;
  assign n225 = ~n220 & ~n224;
  assign n226 = ~\A95  & ~n225;
  assign n227 = ~\A96  & ~n223;
  assign n228 = \A96  & ~n225;
  assign n229 = ~n227 & ~n228;
  assign n230 = \A95  & ~n229;
  assign n231 = ~n226 & ~n230;
  assign n232 = ~\A93  & ~n231;
  assign n233 = ~\A94  & ~n229;
  assign n234 = \A94  & ~n231;
  assign n235 = ~n233 & ~n234;
  assign n236 = \A93  & ~n235;
  assign n237 = ~n232 & ~n236;
  assign n238 = ~\A91  & ~n237;
  assign n239 = ~\A92  & ~n235;
  assign n240 = \A92  & ~n237;
  assign n241 = ~n239 & ~n240;
  assign n242 = \A91  & ~n241;
  assign n243 = ~n238 & ~n242;
  assign n244 = ~\A89  & ~n243;
  assign n245 = ~\A90  & ~n241;
  assign n246 = \A90  & ~n243;
  assign n247 = ~n245 & ~n246;
  assign n248 = \A89  & ~n247;
  assign n249 = ~n244 & ~n248;
  assign n250 = ~\A87  & ~n249;
  assign n251 = ~\A88  & ~n247;
  assign n252 = \A88  & ~n249;
  assign n253 = ~n251 & ~n252;
  assign n254 = \A87  & ~n253;
  assign n255 = ~n250 & ~n254;
  assign n256 = ~\A85  & ~n255;
  assign n257 = ~\A86  & ~n253;
  assign n258 = \A86  & ~n255;
  assign n259 = ~n257 & ~n258;
  assign n260 = \A85  & ~n259;
  assign n261 = ~n256 & ~n260;
  assign n262 = ~\A83  & ~n261;
  assign n263 = ~\A84  & ~n259;
  assign n264 = \A84  & ~n261;
  assign n265 = ~n263 & ~n264;
  assign n266 = \A83  & ~n265;
  assign n267 = ~n262 & ~n266;
  assign n268 = ~\A81  & ~n267;
  assign n269 = ~\A82  & ~n265;
  assign n270 = \A82  & ~n267;
  assign n271 = ~n269 & ~n270;
  assign n272 = \A81  & ~n271;
  assign n273 = ~n268 & ~n272;
  assign n274 = ~\A79  & ~n273;
  assign n275 = ~\A80  & ~n271;
  assign n276 = \A80  & ~n273;
  assign n277 = ~n275 & ~n276;
  assign n278 = \A79  & ~n277;
  assign n279 = ~n274 & ~n278;
  assign n280 = ~\A77  & ~n279;
  assign n281 = ~\A78  & ~n277;
  assign n282 = \A78  & ~n279;
  assign n283 = ~n281 & ~n282;
  assign n284 = \A77  & ~n283;
  assign n285 = ~n280 & ~n284;
  assign n286 = ~\A75  & ~n285;
  assign n287 = ~\A76  & ~n283;
  assign n288 = \A76  & ~n285;
  assign n289 = ~n287 & ~n288;
  assign n290 = \A75  & ~n289;
  assign n291 = ~n286 & ~n290;
  assign n292 = ~\A73  & ~n291;
  assign n293 = ~\A74  & ~n289;
  assign n294 = \A74  & ~n291;
  assign n295 = ~n293 & ~n294;
  assign n296 = \A73  & ~n295;
  assign n297 = ~n292 & ~n296;
  assign n298 = ~\A71  & ~n297;
  assign n299 = ~\A72  & ~n295;
  assign n300 = \A72  & ~n297;
  assign n301 = ~n299 & ~n300;
  assign n302 = \A71  & ~n301;
  assign n303 = ~n298 & ~n302;
  assign n304 = ~\A69  & ~n303;
  assign n305 = ~\A70  & ~n301;
  assign n306 = \A70  & ~n303;
  assign n307 = ~n305 & ~n306;
  assign n308 = \A69  & ~n307;
  assign n309 = ~n304 & ~n308;
  assign n310 = ~\A67  & ~n309;
  assign n311 = ~\A68  & ~n307;
  assign n312 = \A68  & ~n309;
  assign n313 = ~n311 & ~n312;
  assign n314 = \A67  & ~n313;
  assign n315 = ~n310 & ~n314;
  assign n316 = ~\A65  & ~n315;
  assign n317 = ~\A66  & ~n313;
  assign n318 = \A66  & ~n315;
  assign n319 = ~n317 & ~n318;
  assign n320 = \A65  & ~n319;
  assign n321 = ~n316 & ~n320;
  assign n322 = ~\A63  & ~n321;
  assign n323 = ~\A64  & ~n319;
  assign n324 = \A64  & ~n321;
  assign n325 = ~n323 & ~n324;
  assign n326 = \A63  & ~n325;
  assign n327 = ~n322 & ~n326;
  assign n328 = ~\A61  & ~n327;
  assign n329 = ~\A62  & ~n325;
  assign n330 = \A62  & ~n327;
  assign n331 = ~n329 & ~n330;
  assign n332 = \A61  & ~n331;
  assign n333 = ~n328 & ~n332;
  assign n334 = ~\A59  & ~n333;
  assign n335 = ~\A60  & ~n331;
  assign n336 = \A60  & ~n333;
  assign n337 = ~n335 & ~n336;
  assign n338 = \A59  & ~n337;
  assign n339 = ~n334 & ~n338;
  assign n340 = ~\A57  & ~n339;
  assign n341 = ~\A58  & ~n337;
  assign n342 = \A58  & ~n339;
  assign n343 = ~n341 & ~n342;
  assign n344 = \A57  & ~n343;
  assign n345 = ~n340 & ~n344;
  assign n346 = ~\A55  & ~n345;
  assign n347 = ~\A56  & ~n343;
  assign n348 = \A56  & ~n345;
  assign n349 = ~n347 & ~n348;
  assign n350 = \A55  & ~n349;
  assign n351 = ~n346 & ~n350;
  assign n352 = ~\A53  & ~n351;
  assign n353 = ~\A54  & ~n349;
  assign n354 = \A54  & ~n351;
  assign n355 = ~n353 & ~n354;
  assign n356 = \A53  & ~n355;
  assign n357 = ~n352 & ~n356;
  assign n358 = ~\A51  & ~n357;
  assign n359 = ~\A52  & ~n355;
  assign n360 = \A52  & ~n357;
  assign n361 = ~n359 & ~n360;
  assign n362 = \A51  & ~n361;
  assign n363 = ~n358 & ~n362;
  assign n364 = ~\A49  & ~n363;
  assign n365 = ~\A50  & ~n361;
  assign n366 = \A50  & ~n363;
  assign n367 = ~n365 & ~n366;
  assign n368 = \A49  & ~n367;
  assign n369 = ~n364 & ~n368;
  assign n370 = ~\A47  & ~n369;
  assign n371 = ~\A48  & ~n367;
  assign n372 = \A48  & ~n369;
  assign n373 = ~n371 & ~n372;
  assign n374 = \A47  & ~n373;
  assign n375 = ~n370 & ~n374;
  assign n376 = ~\A45  & ~n375;
  assign n377 = ~\A46  & ~n373;
  assign n378 = \A46  & ~n375;
  assign n379 = ~n377 & ~n378;
  assign n380 = \A45  & ~n379;
  assign n381 = ~n376 & ~n380;
  assign n382 = ~\A43  & ~n381;
  assign n383 = ~\A44  & ~n379;
  assign n384 = \A44  & ~n381;
  assign n385 = ~n383 & ~n384;
  assign n386 = \A43  & ~n385;
  assign n387 = ~n382 & ~n386;
  assign n388 = ~\A41  & ~n387;
  assign n389 = ~\A42  & ~n385;
  assign n390 = \A42  & ~n387;
  assign n391 = ~n389 & ~n390;
  assign n392 = \A41  & ~n391;
  assign n393 = ~n388 & ~n392;
  assign n394 = ~\A39  & ~n393;
  assign n395 = ~\A40  & ~n391;
  assign n396 = \A40  & ~n393;
  assign n397 = ~n395 & ~n396;
  assign n398 = \A39  & ~n397;
  assign n399 = ~n394 & ~n398;
  assign n400 = ~\A37  & ~n399;
  assign n401 = ~\A38  & ~n397;
  assign n402 = \A38  & ~n399;
  assign n403 = ~n401 & ~n402;
  assign n404 = \A37  & ~n403;
  assign n405 = ~n400 & ~n404;
  assign n406 = ~\A35  & ~n405;
  assign n407 = ~\A36  & ~n403;
  assign n408 = \A36  & ~n405;
  assign n409 = ~n407 & ~n408;
  assign n410 = \A35  & ~n409;
  assign n411 = ~n406 & ~n410;
  assign n412 = ~\A33  & ~n411;
  assign n413 = ~\A34  & ~n409;
  assign n414 = \A34  & ~n411;
  assign n415 = ~n413 & ~n414;
  assign n416 = \A33  & ~n415;
  assign n417 = ~n412 & ~n416;
  assign n418 = ~\A31  & ~n417;
  assign n419 = ~\A32  & ~n415;
  assign n420 = \A32  & ~n417;
  assign n421 = ~n419 & ~n420;
  assign n422 = \A31  & ~n421;
  assign n423 = ~n418 & ~n422;
  assign n424 = ~\A29  & ~n423;
  assign n425 = ~\A30  & ~n421;
  assign n426 = \A30  & ~n423;
  assign n427 = ~n425 & ~n426;
  assign n428 = \A29  & ~n427;
  assign n429 = ~n424 & ~n428;
  assign n430 = ~\A27  & ~n429;
  assign n431 = ~\A28  & ~n427;
  assign n432 = \A28  & ~n429;
  assign n433 = ~n431 & ~n432;
  assign n434 = \A27  & ~n433;
  assign n435 = ~n430 & ~n434;
  assign n436 = ~\A25  & ~n435;
  assign n437 = ~\A26  & ~n433;
  assign n438 = \A26  & ~n435;
  assign n439 = ~n437 & ~n438;
  assign n440 = \A25  & ~n439;
  assign n441 = ~n436 & ~n440;
  assign n442 = ~\A23  & ~n441;
  assign n443 = ~\A24  & ~n439;
  assign n444 = \A24  & ~n441;
  assign n445 = ~n443 & ~n444;
  assign n446 = \A23  & ~n445;
  assign n447 = ~n442 & ~n446;
  assign n448 = ~\A21  & ~n447;
  assign n449 = ~\A22  & ~n445;
  assign n450 = \A22  & ~n447;
  assign n451 = ~n449 & ~n450;
  assign n452 = \A21  & ~n451;
  assign n453 = ~n448 & ~n452;
  assign n454 = ~\A19  & ~n453;
  assign n455 = ~\A20  & ~n451;
  assign n456 = \A20  & ~n453;
  assign n457 = ~n455 & ~n456;
  assign n458 = \A19  & ~n457;
  assign n459 = ~n454 & ~n458;
  assign n460 = ~\A17  & ~n459;
  assign n461 = ~\A18  & ~n457;
  assign n462 = \A18  & ~n459;
  assign n463 = ~n461 & ~n462;
  assign n464 = \A17  & ~n463;
  assign n465 = ~n460 & ~n464;
  assign n466 = ~\A15  & ~n465;
  assign n467 = ~\A16  & ~n463;
  assign n468 = \A16  & ~n465;
  assign n469 = ~n467 & ~n468;
  assign n470 = \A15  & ~n469;
  assign n471 = ~n466 & ~n470;
  assign n472 = ~\A13  & ~n471;
  assign n473 = ~\A14  & ~n469;
  assign n474 = \A14  & ~n471;
  assign n475 = ~n473 & ~n474;
  assign n476 = \A13  & ~n475;
  assign n477 = ~n472 & ~n476;
  assign n478 = ~\A11  & ~n477;
  assign n479 = ~\A12  & ~n475;
  assign n480 = \A12  & ~n477;
  assign n481 = ~n479 & ~n480;
  assign n482 = \A11  & ~n481;
  assign n483 = ~n478 & ~n482;
  assign n484 = ~\A9  & ~n483;
  assign n485 = ~\A10  & ~n481;
  assign n486 = \A10  & ~n483;
  assign n487 = ~n485 & ~n486;
  assign n488 = \A9  & ~n487;
  assign n489 = ~n484 & ~n488;
  assign n490 = ~\A7  & ~n489;
  assign n491 = ~\A8  & ~n487;
  assign n492 = \A8  & ~n489;
  assign n493 = ~n491 & ~n492;
  assign n494 = \A7  & ~n493;
  assign n495 = ~n490 & ~n494;
  assign n496 = ~\A5  & ~n495;
  assign n497 = ~\A6  & ~n493;
  assign n498 = \A6  & ~n495;
  assign n499 = ~n497 & ~n498;
  assign n500 = \A5  & ~n499;
  assign n501 = ~n496 & ~n500;
  assign n502 = ~\A3  & ~n501;
  assign n503 = ~\A4  & ~n499;
  assign n504 = \A4  & ~n501;
  assign n505 = ~n503 & ~n504;
  assign n506 = \A3  & ~n505;
  assign n507 = ~n502 & ~n506;
  assign n508 = \A1  & ~\A2 ;
  assign n509 = n507 & ~n508;
  assign n510 = n505 & n508;
  assign \P0  = ~n509 & ~n510;
  assign n512 = ~\A126  & \A127 ;
  assign n513 = ~\A126  & ~n512;
  assign n514 = ~\A124  & ~\A125 ;
  assign n515 = ~\A122  & ~\A123 ;
  assign n516 = \A121  & n515;
  assign n517 = n514 & ~n516;
  assign n518 = n513 & ~n517;
  assign n519 = ~\A120  & ~n518;
  assign n520 = n514 & ~n515;
  assign n521 = n513 & ~n520;
  assign n522 = \A120  & ~n521;
  assign n523 = ~n519 & ~n522;
  assign n524 = ~\A118  & ~\A119 ;
  assign n525 = n523 & ~n524;
  assign n526 = n521 & n524;
  assign n527 = ~n525 & ~n526;
  assign n528 = ~\A116  & ~\A117 ;
  assign n529 = n527 & ~n528;
  assign n530 = ~n523 & n528;
  assign n531 = ~n529 & ~n530;
  assign n532 = ~\A114  & ~\A115 ;
  assign n533 = n531 & ~n532;
  assign n534 = ~n527 & n532;
  assign n535 = ~n533 & ~n534;
  assign n536 = ~\A112  & ~\A113 ;
  assign n537 = n535 & ~n536;
  assign n538 = ~n531 & n536;
  assign n539 = ~n537 & ~n538;
  assign n540 = ~\A110  & ~\A111 ;
  assign n541 = n539 & ~n540;
  assign n542 = ~n535 & n540;
  assign n543 = ~n541 & ~n542;
  assign n544 = ~\A108  & ~\A109 ;
  assign n545 = n543 & ~n544;
  assign n546 = ~n539 & n544;
  assign n547 = ~n545 & ~n546;
  assign n548 = ~\A106  & ~\A107 ;
  assign n549 = n547 & ~n548;
  assign n550 = ~n543 & n548;
  assign n551 = ~n549 & ~n550;
  assign n552 = ~\A104  & ~\A105 ;
  assign n553 = n551 & ~n552;
  assign n554 = ~n547 & n552;
  assign n555 = ~n553 & ~n554;
  assign n556 = ~\A102  & ~\A103 ;
  assign n557 = n555 & ~n556;
  assign n558 = ~n551 & n556;
  assign n559 = ~n557 & ~n558;
  assign n560 = ~\A100  & ~\A101 ;
  assign n561 = n559 & ~n560;
  assign n562 = ~n555 & n560;
  assign n563 = ~n561 & ~n562;
  assign n564 = ~\A98  & ~\A99 ;
  assign n565 = n563 & ~n564;
  assign n566 = ~n559 & n564;
  assign n567 = ~n565 & ~n566;
  assign n568 = ~\A96  & ~\A97 ;
  assign n569 = n567 & ~n568;
  assign n570 = ~n563 & n568;
  assign n571 = ~n569 & ~n570;
  assign n572 = ~\A94  & ~\A95 ;
  assign n573 = n571 & ~n572;
  assign n574 = ~n567 & n572;
  assign n575 = ~n573 & ~n574;
  assign n576 = ~\A92  & ~\A93 ;
  assign n577 = n575 & ~n576;
  assign n578 = ~n571 & n576;
  assign n579 = ~n577 & ~n578;
  assign n580 = ~\A90  & ~\A91 ;
  assign n581 = n579 & ~n580;
  assign n582 = ~n575 & n580;
  assign n583 = ~n581 & ~n582;
  assign n584 = ~\A88  & ~\A89 ;
  assign n585 = n583 & ~n584;
  assign n586 = ~n579 & n584;
  assign n587 = ~n585 & ~n586;
  assign n588 = ~\A86  & ~\A87 ;
  assign n589 = n587 & ~n588;
  assign n590 = ~n583 & n588;
  assign n591 = ~n589 & ~n590;
  assign n592 = ~\A84  & ~\A85 ;
  assign n593 = n591 & ~n592;
  assign n594 = ~n587 & n592;
  assign n595 = ~n593 & ~n594;
  assign n596 = ~\A82  & ~\A83 ;
  assign n597 = n595 & ~n596;
  assign n598 = ~n591 & n596;
  assign n599 = ~n597 & ~n598;
  assign n600 = ~\A80  & ~\A81 ;
  assign n601 = n599 & ~n600;
  assign n602 = ~n595 & n600;
  assign n603 = ~n601 & ~n602;
  assign n604 = ~\A78  & ~\A79 ;
  assign n605 = n603 & ~n604;
  assign n606 = ~n599 & n604;
  assign n607 = ~n605 & ~n606;
  assign n608 = ~\A76  & ~\A77 ;
  assign n609 = n607 & ~n608;
  assign n610 = ~n603 & n608;
  assign n611 = ~n609 & ~n610;
  assign n612 = ~\A74  & ~\A75 ;
  assign n613 = n611 & ~n612;
  assign n614 = ~n607 & n612;
  assign n615 = ~n613 & ~n614;
  assign n616 = ~\A72  & ~\A73 ;
  assign n617 = n615 & ~n616;
  assign n618 = ~n611 & n616;
  assign n619 = ~n617 & ~n618;
  assign n620 = ~\A70  & ~\A71 ;
  assign n621 = n619 & ~n620;
  assign n622 = ~n615 & n620;
  assign n623 = ~n621 & ~n622;
  assign n624 = ~\A68  & ~\A69 ;
  assign n625 = n623 & ~n624;
  assign n626 = ~n619 & n624;
  assign n627 = ~n625 & ~n626;
  assign n628 = ~\A66  & ~\A67 ;
  assign n629 = n627 & ~n628;
  assign n630 = ~n623 & n628;
  assign n631 = ~n629 & ~n630;
  assign n632 = ~\A64  & ~\A65 ;
  assign n633 = n631 & ~n632;
  assign n634 = ~n627 & n632;
  assign n635 = ~n633 & ~n634;
  assign n636 = ~\A62  & ~\A63 ;
  assign n637 = n635 & ~n636;
  assign n638 = ~n631 & n636;
  assign n639 = ~n637 & ~n638;
  assign n640 = ~\A60  & ~\A61 ;
  assign n641 = n639 & ~n640;
  assign n642 = ~n635 & n640;
  assign n643 = ~n641 & ~n642;
  assign n644 = ~\A58  & ~\A59 ;
  assign n645 = n643 & ~n644;
  assign n646 = ~n639 & n644;
  assign n647 = ~n645 & ~n646;
  assign n648 = ~\A56  & ~\A57 ;
  assign n649 = n647 & ~n648;
  assign n650 = ~n643 & n648;
  assign n651 = ~n649 & ~n650;
  assign n652 = ~\A54  & ~\A55 ;
  assign n653 = n651 & ~n652;
  assign n654 = ~n647 & n652;
  assign n655 = ~n653 & ~n654;
  assign n656 = ~\A52  & ~\A53 ;
  assign n657 = n655 & ~n656;
  assign n658 = ~n651 & n656;
  assign n659 = ~n657 & ~n658;
  assign n660 = ~\A50  & ~\A51 ;
  assign n661 = n659 & ~n660;
  assign n662 = ~n655 & n660;
  assign n663 = ~n661 & ~n662;
  assign n664 = ~\A48  & ~\A49 ;
  assign n665 = n663 & ~n664;
  assign n666 = ~n659 & n664;
  assign n667 = ~n665 & ~n666;
  assign n668 = ~\A46  & ~\A47 ;
  assign n669 = n667 & ~n668;
  assign n670 = ~n663 & n668;
  assign n671 = ~n669 & ~n670;
  assign n672 = ~\A44  & ~\A45 ;
  assign n673 = n671 & ~n672;
  assign n674 = ~n667 & n672;
  assign n675 = ~n673 & ~n674;
  assign n676 = ~\A42  & ~\A43 ;
  assign n677 = n675 & ~n676;
  assign n678 = ~n671 & n676;
  assign n679 = ~n677 & ~n678;
  assign n680 = ~\A40  & ~\A41 ;
  assign n681 = n679 & ~n680;
  assign n682 = ~n675 & n680;
  assign n683 = ~n681 & ~n682;
  assign n684 = ~\A38  & ~\A39 ;
  assign n685 = n683 & ~n684;
  assign n686 = ~n679 & n684;
  assign n687 = ~n685 & ~n686;
  assign n688 = ~\A36  & ~\A37 ;
  assign n689 = n687 & ~n688;
  assign n690 = ~n683 & n688;
  assign n691 = ~n689 & ~n690;
  assign n692 = ~\A34  & ~\A35 ;
  assign n693 = n691 & ~n692;
  assign n694 = ~n687 & n692;
  assign n695 = ~n693 & ~n694;
  assign n696 = ~\A32  & ~\A33 ;
  assign n697 = n695 & ~n696;
  assign n698 = ~n691 & n696;
  assign n699 = ~n697 & ~n698;
  assign n700 = ~\A30  & ~\A31 ;
  assign n701 = n699 & ~n700;
  assign n702 = ~n695 & n700;
  assign n703 = ~n701 & ~n702;
  assign n704 = ~\A28  & ~\A29 ;
  assign n705 = n703 & ~n704;
  assign n706 = ~n699 & n704;
  assign n707 = ~n705 & ~n706;
  assign n708 = ~\A26  & ~\A27 ;
  assign n709 = n707 & ~n708;
  assign n710 = ~n703 & n708;
  assign n711 = ~n709 & ~n710;
  assign n712 = ~\A24  & ~\A25 ;
  assign n713 = n711 & ~n712;
  assign n714 = ~n707 & n712;
  assign n715 = ~n713 & ~n714;
  assign n716 = ~\A22  & ~\A23 ;
  assign n717 = n715 & ~n716;
  assign n718 = ~n711 & n716;
  assign n719 = ~n717 & ~n718;
  assign n720 = ~\A20  & ~\A21 ;
  assign n721 = n719 & ~n720;
  assign n722 = ~n715 & n720;
  assign n723 = ~n721 & ~n722;
  assign n724 = ~\A18  & ~\A19 ;
  assign n725 = n723 & ~n724;
  assign n726 = ~n719 & n724;
  assign n727 = ~n725 & ~n726;
  assign n728 = ~\A16  & ~\A17 ;
  assign n729 = n727 & ~n728;
  assign n730 = ~n723 & n728;
  assign n731 = ~n729 & ~n730;
  assign n732 = ~\A14  & ~\A15 ;
  assign n733 = n731 & ~n732;
  assign n734 = ~n727 & n732;
  assign n735 = ~n733 & ~n734;
  assign n736 = ~\A12  & ~\A13 ;
  assign n737 = n735 & ~n736;
  assign n738 = ~n731 & n736;
  assign n739 = ~n737 & ~n738;
  assign n740 = ~\A10  & ~\A11 ;
  assign n741 = n739 & ~n740;
  assign n742 = ~n735 & n740;
  assign n743 = ~n741 & ~n742;
  assign n744 = ~\A8  & ~\A9 ;
  assign n745 = n743 & ~n744;
  assign n746 = ~n739 & n744;
  assign n747 = ~n745 & ~n746;
  assign n748 = ~\A6  & ~\A7 ;
  assign n749 = n747 & ~n748;
  assign n750 = ~n743 & n748;
  assign n751 = ~n749 & ~n750;
  assign n752 = ~\A4  & ~\A5 ;
  assign n753 = n751 & ~n752;
  assign n754 = ~n747 & n752;
  assign n755 = ~n753 & ~n754;
  assign n756 = ~\A2  & ~\A3 ;
  assign n757 = n755 & ~n756;
  assign n758 = ~n751 & n756;
  assign \P1  = ~n757 & ~n758;
  assign n760 = n513 & n514;
  assign n761 = ~\A120  & ~\A121 ;
  assign n762 = n515 & n761;
  assign n763 = ~\A117  & n524;
  assign n764 = ~\A116  & n763;
  assign n765 = n762 & ~n764;
  assign n766 = n760 & ~n765;
  assign n767 = ~\A113  & ~\A114 ;
  assign n768 = ~\A112  & n767;
  assign n769 = n766 & ~n768;
  assign n770 = \A115  & n764;
  assign n771 = n762 & ~n770;
  assign n772 = n760 & ~n771;
  assign n773 = n768 & n772;
  assign n774 = ~n769 & ~n773;
  assign n775 = ~\A109  & n540;
  assign n776 = ~\A108  & n775;
  assign n777 = n774 & ~n776;
  assign n778 = ~n766 & n776;
  assign n779 = ~n777 & ~n778;
  assign n780 = ~\A105  & n548;
  assign n781 = ~\A104  & n780;
  assign n782 = n779 & ~n781;
  assign n783 = ~n774 & n781;
  assign n784 = ~n782 & ~n783;
  assign n785 = ~\A101  & n556;
  assign n786 = ~\A100  & n785;
  assign n787 = n784 & ~n786;
  assign n788 = ~n779 & n786;
  assign n789 = ~n787 & ~n788;
  assign n790 = ~\A97  & n564;
  assign n791 = ~\A96  & n790;
  assign n792 = n789 & ~n791;
  assign n793 = ~n784 & n791;
  assign n794 = ~n792 & ~n793;
  assign n795 = ~\A93  & n572;
  assign n796 = ~\A92  & n795;
  assign n797 = n794 & ~n796;
  assign n798 = ~n789 & n796;
  assign n799 = ~n797 & ~n798;
  assign n800 = ~\A89  & n580;
  assign n801 = ~\A88  & n800;
  assign n802 = n799 & ~n801;
  assign n803 = ~n794 & n801;
  assign n804 = ~n802 & ~n803;
  assign n805 = ~\A85  & n588;
  assign n806 = ~\A84  & n805;
  assign n807 = n804 & ~n806;
  assign n808 = ~n799 & n806;
  assign n809 = ~n807 & ~n808;
  assign n810 = ~\A81  & n596;
  assign n811 = ~\A80  & n810;
  assign n812 = n809 & ~n811;
  assign n813 = ~n804 & n811;
  assign n814 = ~n812 & ~n813;
  assign n815 = ~\A77  & n604;
  assign n816 = ~\A76  & n815;
  assign n817 = n814 & ~n816;
  assign n818 = ~n809 & n816;
  assign n819 = ~n817 & ~n818;
  assign n820 = ~\A73  & n612;
  assign n821 = ~\A72  & n820;
  assign n822 = n819 & ~n821;
  assign n823 = ~n814 & n821;
  assign n824 = ~n822 & ~n823;
  assign n825 = ~\A69  & n620;
  assign n826 = ~\A68  & n825;
  assign n827 = n824 & ~n826;
  assign n828 = ~n819 & n826;
  assign n829 = ~n827 & ~n828;
  assign n830 = ~\A65  & n628;
  assign n831 = ~\A64  & n830;
  assign n832 = n829 & ~n831;
  assign n833 = ~n824 & n831;
  assign n834 = ~n832 & ~n833;
  assign n835 = ~\A61  & n636;
  assign n836 = ~\A60  & n835;
  assign n837 = n834 & ~n836;
  assign n838 = ~n829 & n836;
  assign n839 = ~n837 & ~n838;
  assign n840 = ~\A57  & n644;
  assign n841 = ~\A56  & n840;
  assign n842 = n839 & ~n841;
  assign n843 = ~n834 & n841;
  assign n844 = ~n842 & ~n843;
  assign n845 = ~\A53  & n652;
  assign n846 = ~\A52  & n845;
  assign n847 = n844 & ~n846;
  assign n848 = ~n839 & n846;
  assign n849 = ~n847 & ~n848;
  assign n850 = ~\A49  & n660;
  assign n851 = ~\A48  & n850;
  assign n852 = n849 & ~n851;
  assign n853 = ~n844 & n851;
  assign n854 = ~n852 & ~n853;
  assign n855 = ~\A45  & n668;
  assign n856 = ~\A44  & n855;
  assign n857 = n854 & ~n856;
  assign n858 = ~n849 & n856;
  assign n859 = ~n857 & ~n858;
  assign n860 = ~\A41  & n676;
  assign n861 = ~\A40  & n860;
  assign n862 = n859 & ~n861;
  assign n863 = ~n854 & n861;
  assign n864 = ~n862 & ~n863;
  assign n865 = ~\A37  & n684;
  assign n866 = ~\A36  & n865;
  assign n867 = n864 & ~n866;
  assign n868 = ~n859 & n866;
  assign n869 = ~n867 & ~n868;
  assign n870 = ~\A33  & n692;
  assign n871 = ~\A32  & n870;
  assign n872 = n869 & ~n871;
  assign n873 = ~n864 & n871;
  assign n874 = ~n872 & ~n873;
  assign n875 = ~\A29  & n700;
  assign n876 = ~\A28  & n875;
  assign n877 = n874 & ~n876;
  assign n878 = ~n869 & n876;
  assign n879 = ~n877 & ~n878;
  assign n880 = ~\A25  & n708;
  assign n881 = ~\A24  & n880;
  assign n882 = n879 & ~n881;
  assign n883 = ~n874 & n881;
  assign n884 = ~n882 & ~n883;
  assign n885 = ~\A21  & n716;
  assign n886 = ~\A20  & n885;
  assign n887 = n884 & ~n886;
  assign n888 = ~n879 & n886;
  assign n889 = ~n887 & ~n888;
  assign n890 = ~\A17  & n724;
  assign n891 = ~\A16  & n890;
  assign n892 = n889 & ~n891;
  assign n893 = ~n884 & n891;
  assign n894 = ~n892 & ~n893;
  assign n895 = ~\A13  & n732;
  assign n896 = ~\A12  & n895;
  assign n897 = n894 & ~n896;
  assign n898 = ~n889 & n896;
  assign n899 = ~n897 & ~n898;
  assign n900 = ~\A9  & n740;
  assign n901 = ~\A8  & n900;
  assign n902 = n899 & ~n901;
  assign n903 = ~n894 & n901;
  assign n904 = ~n902 & ~n903;
  assign n905 = ~\A5  & n748;
  assign n906 = ~\A4  & n905;
  assign n907 = n904 & ~n906;
  assign n908 = ~n899 & n906;
  assign \P2  = n907 | n908;
  assign n910 = n760 & n762;
  assign n911 = ~\A113  & n532;
  assign n912 = ~\A112  & n764;
  assign n913 = n911 & n912;
  assign n914 = ~\A107  & n776;
  assign n915 = ~\A106  & n914;
  assign n916 = ~\A105  & n915;
  assign n917 = ~\A104  & n916;
  assign n918 = n913 & ~n917;
  assign n919 = n910 & ~n918;
  assign n920 = ~\A101  & ~\A102 ;
  assign n921 = ~\A100  & n920;
  assign n922 = ~\A99  & n921;
  assign n923 = ~\A98  & n922;
  assign n924 = ~\A97  & n923;
  assign n925 = ~\A96  & n924;
  assign n926 = n919 & ~n925;
  assign n927 = \A103  & n917;
  assign n928 = n913 & ~n927;
  assign n929 = n910 & ~n928;
  assign n930 = n925 & n929;
  assign n931 = ~n926 & ~n930;
  assign n932 = ~\A91  & n796;
  assign n933 = ~\A90  & n932;
  assign n934 = ~\A89  & n933;
  assign n935 = ~\A88  & n934;
  assign n936 = n931 & ~n935;
  assign n937 = ~n919 & n935;
  assign n938 = ~n936 & ~n937;
  assign n939 = ~\A83  & n806;
  assign n940 = ~\A82  & n939;
  assign n941 = ~\A81  & n940;
  assign n942 = ~\A80  & n941;
  assign n943 = n938 & ~n942;
  assign n944 = ~n931 & n942;
  assign n945 = ~n943 & ~n944;
  assign n946 = ~\A75  & n816;
  assign n947 = ~\A74  & n946;
  assign n948 = ~\A73  & n947;
  assign n949 = ~\A72  & n948;
  assign n950 = n945 & ~n949;
  assign n951 = ~n938 & n949;
  assign n952 = ~n950 & ~n951;
  assign n953 = ~\A67  & n826;
  assign n954 = ~\A66  & n953;
  assign n955 = ~\A65  & n954;
  assign n956 = ~\A64  & n955;
  assign n957 = n952 & ~n956;
  assign n958 = ~n945 & n956;
  assign n959 = ~n957 & ~n958;
  assign n960 = ~\A59  & n836;
  assign n961 = ~\A58  & n960;
  assign n962 = ~\A57  & n961;
  assign n963 = ~\A56  & n962;
  assign n964 = n959 & ~n963;
  assign n965 = ~n952 & n963;
  assign n966 = ~n964 & ~n965;
  assign n967 = ~\A51  & n846;
  assign n968 = ~\A50  & n967;
  assign n969 = ~\A49  & n968;
  assign n970 = ~\A48  & n969;
  assign n971 = n966 & ~n970;
  assign n972 = ~n959 & n970;
  assign n973 = ~n971 & ~n972;
  assign n974 = ~\A43  & n856;
  assign n975 = ~\A42  & n974;
  assign n976 = ~\A41  & n975;
  assign n977 = ~\A40  & n976;
  assign n978 = n973 & ~n977;
  assign n979 = ~n966 & n977;
  assign n980 = ~n978 & ~n979;
  assign n981 = ~\A35  & n866;
  assign n982 = ~\A34  & n981;
  assign n983 = ~\A33  & n982;
  assign n984 = ~\A32  & n983;
  assign n985 = n980 & ~n984;
  assign n986 = ~n973 & n984;
  assign n987 = ~n985 & ~n986;
  assign n988 = ~\A27  & n876;
  assign n989 = ~\A26  & n988;
  assign n990 = ~\A25  & n989;
  assign n991 = ~\A24  & n990;
  assign n992 = n987 & ~n991;
  assign n993 = ~n980 & n991;
  assign n994 = ~n992 & ~n993;
  assign n995 = ~\A19  & n886;
  assign n996 = ~\A18  & n995;
  assign n997 = ~\A17  & n996;
  assign n998 = ~\A16  & n997;
  assign n999 = n994 & ~n998;
  assign n1000 = ~n987 & n998;
  assign n1001 = ~n999 & ~n1000;
  assign n1002 = ~\A11  & n896;
  assign n1003 = ~\A10  & n1002;
  assign n1004 = ~\A9  & n1003;
  assign n1005 = ~\A8  & n1004;
  assign n1006 = n1001 & ~n1005;
  assign n1007 = ~n994 & n1005;
  assign \P3  = n1006 | n1007;
  assign n1009 = n910 & n913;
  assign n1010 = ~\A99  & n786;
  assign n1011 = ~\A98  & n917;
  assign n1012 = ~\A97  & n1011;
  assign n1013 = ~\A96  & n1012;
  assign n1014 = n1010 & n1013;
  assign n1015 = ~\A87  & n935;
  assign n1016 = ~\A86  & n1015;
  assign n1017 = ~\A85  & n1016;
  assign n1018 = ~\A84  & n1017;
  assign n1019 = ~\A83  & n1018;
  assign n1020 = ~\A82  & n1019;
  assign n1021 = ~\A81  & n1020;
  assign n1022 = ~\A80  & n1021;
  assign n1023 = n1014 & ~n1022;
  assign n1024 = n1009 & ~n1023;
  assign n1025 = ~\A77  & ~\A78 ;
  assign n1026 = ~\A76  & n1025;
  assign n1027 = ~\A75  & n1026;
  assign n1028 = ~\A74  & n1027;
  assign n1029 = ~\A73  & n1028;
  assign n1030 = ~\A72  & n1029;
  assign n1031 = ~\A71  & n1030;
  assign n1032 = ~\A70  & n1031;
  assign n1033 = ~\A69  & n1032;
  assign n1034 = ~\A68  & n1033;
  assign n1035 = ~\A67  & n1034;
  assign n1036 = ~\A66  & n1035;
  assign n1037 = ~\A65  & n1036;
  assign n1038 = ~\A64  & n1037;
  assign n1039 = n1024 & ~n1038;
  assign n1040 = \A79  & n1022;
  assign n1041 = n1014 & ~n1040;
  assign n1042 = n1009 & ~n1041;
  assign n1043 = n1038 & n1042;
  assign n1044 = ~n1039 & ~n1043;
  assign n1045 = ~\A55  & n963;
  assign n1046 = ~\A54  & n1045;
  assign n1047 = ~\A53  & n1046;
  assign n1048 = ~\A52  & n1047;
  assign n1049 = ~\A51  & n1048;
  assign n1050 = ~\A50  & n1049;
  assign n1051 = ~\A49  & n1050;
  assign n1052 = ~\A48  & n1051;
  assign n1053 = n1044 & ~n1052;
  assign n1054 = ~n1024 & n1052;
  assign n1055 = ~n1053 & ~n1054;
  assign n1056 = ~\A39  & n977;
  assign n1057 = ~\A38  & n1056;
  assign n1058 = ~\A37  & n1057;
  assign n1059 = ~\A36  & n1058;
  assign n1060 = ~\A35  & n1059;
  assign n1061 = ~\A34  & n1060;
  assign n1062 = ~\A33  & n1061;
  assign n1063 = ~\A32  & n1062;
  assign n1064 = n1055 & ~n1063;
  assign n1065 = ~n1044 & n1063;
  assign n1066 = ~n1064 & ~n1065;
  assign n1067 = ~\A23  & n991;
  assign n1068 = ~\A22  & n1067;
  assign n1069 = ~\A21  & n1068;
  assign n1070 = ~\A20  & n1069;
  assign n1071 = ~\A19  & n1070;
  assign n1072 = ~\A18  & n1071;
  assign n1073 = ~\A17  & n1072;
  assign n1074 = ~\A16  & n1073;
  assign n1075 = n1066 & ~n1074;
  assign n1076 = ~n1055 & n1074;
  assign \P4  = n1075 | n1076;
  assign n1078 = n1009 & n1014;
  assign n1079 = ~\A71  & n949;
  assign n1080 = ~\A70  & n1022;
  assign n1081 = ~\A69  & n1080;
  assign n1082 = ~\A68  & n1081;
  assign n1083 = ~\A67  & n1082;
  assign n1084 = ~\A66  & n1083;
  assign n1085 = ~\A65  & n1084;
  assign n1086 = ~\A64  & n1085;
  assign n1087 = n1079 & n1086;
  assign n1088 = ~\A47  & n1052;
  assign n1089 = ~\A46  & n1088;
  assign n1090 = ~\A45  & n1089;
  assign n1091 = ~\A44  & n1090;
  assign n1092 = ~\A43  & n1091;
  assign n1093 = ~\A42  & n1092;
  assign n1094 = ~\A41  & n1093;
  assign n1095 = ~\A40  & n1094;
  assign n1096 = ~\A39  & n1095;
  assign n1097 = ~\A38  & n1096;
  assign n1098 = ~\A37  & n1097;
  assign n1099 = ~\A36  & n1098;
  assign n1100 = ~\A35  & n1099;
  assign n1101 = ~\A34  & n1100;
  assign n1102 = ~\A33  & n1101;
  assign n1103 = ~\A32  & n1102;
  assign n1104 = n1087 & ~n1103;
  assign \P5  = ~n1078 | n1104;
  assign \P6  = ~n1078 | ~n1087;
  assign n1107 = ~\A0  & ~\P6 ;
  assign n1108 = n1005 & n1107;
  assign n1109 = ~\A3  & n1108;
  assign n1110 = ~\A2  & n1109;
  assign n1111 = n1074 & n1103;
  assign n1112 = n906 & n1111;
  assign n1113 = ~\A1  & n1112;
  assign F = ~n1110 | ~n1113;
endmodule
