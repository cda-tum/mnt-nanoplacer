module top (
    \1 , 4, 11, 14, 17, 20, 23, 24, 25, 26, 27, 31, 34, 37, 40, 43, 46, 49,
    52, 53, 54, 61, 64, 67, 70, 73, 76, 79, 80, 81, 82, 83, 86, 87, 88, 91,
    94, 97, 100, 103, 106, 109, 112, 113, 114, 115, 116, 117, 118, 119,
    120, 121, 122, 123, 126, 127, 128, 129, 130, 131, 132, 135, 136, 137,
    140, 141, 145, 146, 149, 152, 155, 158, 161, 164, 167, 170, 173, 176,
    179, 182, 185, 188, 191, 194, 197, 200, 203, 206, 209, 210, 217, 218,
    225, 226, 233, 234, 241, 242, 245, 248, 251, 254, 257, 264, 265, 272,
    273, 280, 281, 288, 289, 292, 293, 299, 302, 307, 308, 315, 316, 323,
    324, 331, 332, 335, 338, 341, 348, 351, 358, 361, 366, 369, 372, 373,
    374, 386, 389, 400, 411, 422, 435, 446, 457, 468, 479, 490, 503, 514,
    523, 534, 545, 549, 552, 556, 559, 562, 566, 571, 574, 577, 580, 583,
    588, 591, 592, 595, 596, 597, 598, 599, 603, 607, 610, 613, 616, 619,
    625, 631,
    709, 816, 1066, 1137, 1138, 1139, 1140, 1141, 1142, 1143, 1144, 1145,
    1147, 1152, 1153, 1154, 1155, 1972, 2054, 2060, 2061, 2139, 2142, 2309,
    2387, 2527, 2584, 2590, 2623, 3357, 3358, 3359, 3360, 3604, 3613, 4272,
    4275, 4278, 4279, 4737, 4738, 4739, 4740, 5240, 5388, 6641, 6643, 6646,
    6648, 6716, 6877, 6924, 6925, 6926, 6927, 7015, 7363, 7365, 7432, 7449,
    7465, 7466, 7467, 7469, 7470, 7471, 7472, 7473, 7474, 7476, 7503, 7504,
    7506, 7511, 7515, 7516, 7517, 7518, 7519, 7520, 7521, 7522, 7600, 7601,
    7602, 7603, 7604, 7605, 7606, 7607, 7626, 7698, 7699, 7700, 7701, 7702,
    7703, 7704, 7705, 7706, 7707, 7735, 7736, 7737, 7738, 7739, 7740, 7741,
    7742, 7754, 7755, 7756, 7757, 7758, 7759, 7760, 7761, 8075, 8076, 8123,
    8124, 8127, 8128  );
  input  \1 , 4, 11, 14, 17, 20, 23, 24, 25, 26, 27, 31, 34, 37, 40, 43,
    46, 49, 52, 53, 54, 61, 64, 67, 70, 73, 76, 79, 80, 81, 82, 83, 86, 87,
    88, 91, 94, 97, 100, 103, 106, 109, 112, 113, 114, 115, 116, 117, 118,
    119, 120, 121, 122, 123, 126, 127, 128, 129, 130, 131, 132, 135, 136,
    137, 140, 141, 145, 146, 149, 152, 155, 158, 161, 164, 167, 170, 173,
    176, 179, 182, 185, 188, 191, 194, 197, 200, 203, 206, 209, 210, 217,
    218, 225, 226, 233, 234, 241, 242, 245, 248, 251, 254, 257, 264, 265,
    272, 273, 280, 281, 288, 289, 292, 293, 299, 302, 307, 308, 315, 316,
    323, 324, 331, 332, 335, 338, 341, 348, 351, 358, 361, 366, 369, 372,
    373, 374, 386, 389, 400, 411, 422, 435, 446, 457, 468, 479, 490, 503,
    514, 523, 534, 545, 549, 552, 556, 559, 562, 566, 571, 574, 577, 580,
    583, 588, 591, 592, 595, 596, 597, 598, 599, 603, 607, 610, 613, 616,
    619, 625, 631;
  output 709, 816, 1066, 1137, 1138, 1139, 1140, 1141, 1142, 1143, 1144, 1145,
    1147, 1152, 1153, 1154, 1155, 1972, 2054, 2060, 2061, 2139, 2142, 2309,
    2387, 2527, 2584, 2590, 2623, 3357, 3358, 3359, 3360, 3604, 3613, 4272,
    4275, 4278, 4279, 4737, 4738, 4739, 4740, 5240, 5388, 6641, 6643, 6646,
    6648, 6716, 6877, 6924, 6925, 6926, 6927, 7015, 7363, 7365, 7432, 7449,
    7465, 7466, 7467, 7469, 7470, 7471, 7472, 7473, 7474, 7476, 7503, 7504,
    7506, 7511, 7515, 7516, 7517, 7518, 7519, 7520, 7521, 7522, 7600, 7601,
    7602, 7603, 7604, 7605, 7606, 7607, 7626, 7698, 7699, 7700, 7701, 7702,
    7703, 7704, 7705, 7706, 7707, 7735, 7736, 7737, 7738, 7739, 7740, 7741,
    7742, 7754, 7755, 7756, 7757, 7758, 7759, 7760, 7761, 8075, 8076, 8123,
    8124, 8127, 8128;
  wire n310, n311, n312, n314, n315, n316, n318, n319, n320, n322, n323,
    n324, n325, n326, n327, n328, n329, n330, n332, n333, n334, n335, n336,
    n337, n338, n340, n341, n342, n343, n344, n345, n346, n348, n349, n350,
    n351, n352, n353, n354, n356, n357, n358, n359, n360, n361, n362, n363,
    n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
    n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
    n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
    n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
    n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
    n424, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
    n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
    n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
    n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
    n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
    n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
    n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
    n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
    n521, n522, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
    n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
    n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
    n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
    n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
    n582, n583, n584, n586, n587, n588, n589, n590, n591, n592, n593, n594,
    n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
    n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
    n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
    n631, n632, n633, n634, n635, n636, n638, n639, n640, n641, n642, n643,
    n644, n646, n647, n648, n649, n650, n651, n652, n654, n655, n656, n657,
    n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
    n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
    n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
    n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
    n707, n708, n709, n710, n711, n712, n713, n715, n716, n717, n718, n719,
    n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
    n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
    n744, n745, n746, n747, n749, n750, n751, n752, n753, n754, n755, n756,
    n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
    n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n780, n782,
    n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n795, n796,
    n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n808, n809,
    n810, n811, n812, n813, n814, n815, n816, n817, n819, n820, n821, n822,
    n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
    n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n847, n848,
    n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
    n861, n862, n863, n864, n865, n866, n867, n868, n870, n871, n872, n873,
    n874, n875, n876, n877, n878, n879, n880, n881, n882, n884, n885, n886,
    n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n899,
    n900, n901, n902, n903, n904, n905, n906, n907, n908, n910, n911, n912,
    n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924,
    n925, n926, n927, n928, n929, n930, n931, n932, n934, n935, n936, n937,
    n938, n939, n940, n941, n942, n943, n944, n945, n946, n948, n949, n950,
    n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n963,
    n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n975, n976,
    n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988,
    n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999,
    n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1009, n1010,
    n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020,
    n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030,
    n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040,
    n1041, n1042, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051,
    n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061,
    n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071,
    n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081,
    n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091,
    n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
    n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
    n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
    n1123, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
    n1134, n1135, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
    n1145, n1146, n1147, n1149, n1150, n1151, n1152, n1153, n1154, n1155,
    n1156, n1157, n1158, n1160, n1161, n1162, n1163, n1164, n1165, n1166,
    n1167, n1168, n1169, n1171, n1172, n1173, n1174, n1175, n1176, n1177,
    n1178, n1179, n1180, n1182, n1183, n1184, n1185, n1186, n1187, n1188,
    n1189, n1190, n1191, n1193, n1194, n1195, n1196, n1197, n1198, n1199,
    n1200, n1201, n1202, n1204, n1205, n1206, n1207, n1208, n1209, n1210,
    n1211, n1212, n1213, n1215, n1216, n1217, n1218, n1219, n1220, n1221,
    n1222, n1223, n1224, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
    n1233, n1234, n1235, n1237, n1238, n1239, n1240, n1241, n1242, n1243,
    n1244, n1245, n1246, n1247, n1249, n1250, n1251, n1252, n1253, n1254,
    n1255, n1256, n1257, n1258, n1259, n1261, n1262, n1263, n1264, n1265,
    n1266, n1267, n1268, n1269, n1270, n1271, n1273, n1274, n1275, n1276,
    n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1285, n1286, n1287,
    n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1297, n1298,
    n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1309,
    n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319,
    n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330,
    n1331, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341,
    n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1350, n1351, n1352,
    n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1362, n1363, n1364,
    n1365, n1366, n1367, n1368, n1370, n1371, n1372, n1373, n1374, n1375,
    n1376, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1386, n1387,
    n1388, n1389, n1390, n1391, n1392, n1393, n1395, n1396, n1397, n1398,
    n1399, n1400, n1401, n1403, n1404, n1405, n1406, n1407, n1408, n1409,
    n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1419, n1420, n1421,
    n1422, n1423, n1424, n1425, n1427, n1428, n1429, n1430, n1431, n1432,
    n1433, n1434, n1435, n1436, n1438, n1439, n1440, n1441, n1442, n1443,
    n1444, n1445, n1446, n1447, n1449, n1450, n1451, n1452, n1453, n1454,
    n1455, n1456, n1457, n1458, n1460, n1461, n1462, n1463, n1464, n1465,
    n1466, n1467, n1468, n1469, n1471, n1472, n1473, n1474, n1475, n1476,
    n1477, n1478, n1479, n1480, n1482, n1483, n1484, n1485, n1486, n1487,
    n1488, n1489, n1490, n1491, n1493, n1494, n1495, n1496, n1497, n1498,
    n1499, n1500, n1501, n1502, n1504, n1505, n1506, n1507, n1508, n1509,
    n1510, n1511, n1512, n1513, n1515, n1516, n1517, n1518, n1519, n1520,
    n1521, n1522, n1523, n1524, n1525, n1527, n1528, n1529, n1530, n1531,
    n1532, n1533, n1534, n1535, n1536, n1537, n1539, n1540, n1541, n1542,
    n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1551, n1552, n1553,
    n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1563, n1564,
    n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1575,
    n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585,
    n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596,
    n1597, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607,
    n1608, n1609, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618,
    n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628,
    n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638,
    n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648,
    n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658,
    n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668,
    n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678,
    n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688,
    n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698,
    n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708,
    n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718,
    n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728,
    n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738,
    n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748,
    n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758,
    n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768,
    n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778,
    n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1789,
    n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799,
    n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809,
    n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819,
    n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829,
    n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839,
    n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849,
    n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859,
    n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869,
    n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879,
    n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889,
    n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899,
    n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909,
    n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919,
    n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929,
    n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939,
    n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949,
    n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959,
    n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969,
    n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979,
    n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989,
    n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999,
    n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009,
    n2010, n2011, n2012, n2013, n2014, n2015, n2017, n2018, n2019, n2020,
    n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030,
    n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2040, n2041,
    n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2051, n2052,
    n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2063,
    n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073;
  assign 1140 = 552 & 562;
  assign 1147 = 141 & 145;
  assign 1972 = \1  & 373;
  assign 2054 = 136 & ~592;
  assign 2060 = ~27 | 591;
  assign 2061 = ~386 | ~556;
  assign 2623 = ~27 | ~31;
  assign 2590 = ~140 | 2623;
  assign n310 = 87 & 588;
  assign n311 = 86 & ~588;
  assign n312 = ~n310 & ~n311;
  assign 4272 = 2623 | n312;
  assign n314 = 34 & 588;
  assign n315 = 88 & ~588;
  assign n316 = ~n314 & ~n315;
  assign 4275 = 2623 | n316;
  assign n318 = 83 & 588;
  assign n319 = 83 & ~588;
  assign n320 = ~n318 & ~n319;
  assign 4279 = 2623 | n320;
  assign n322 = 24 & ~588;
  assign n323 = ~2623 & n322;
  assign n324 = 25 & 588;
  assign n325 = ~2623 & n324;
  assign n326 = ~588 & 2623;
  assign n327 = 588 & 2623;
  assign n328 = ~n323 & ~n325;
  assign n329 = ~n326 & n328;
  assign n330 = ~n327 & n329;
  assign 4737 = 141 & ~n330;
  assign n332 = 26 & ~588;
  assign n333 = ~2623 & n332;
  assign n334 = 81 & 588;
  assign n335 = ~2623 & n334;
  assign n336 = ~n333 & ~n335;
  assign n337 = ~n326 & n336;
  assign n338 = ~n327 & n337;
  assign 4738 = 141 & ~n338;
  assign n340 = 79 & ~588;
  assign n341 = ~2623 & n340;
  assign n342 = 23 & 588;
  assign n343 = ~2623 & n342;
  assign n344 = ~n341 & ~n343;
  assign n345 = ~n326 & n344;
  assign n346 = ~n327 & n345;
  assign 4739 = 141 & ~n346;
  assign n348 = 82 & ~588;
  assign n349 = ~2623 & n348;
  assign n350 = 80 & 588;
  assign n351 = ~2623 & n350;
  assign n352 = ~n349 & ~n351;
  assign n353 = ~n326 & n352;
  assign n354 = ~n327 & n353;
  assign 4740 = 141 & ~n354;
  assign n356 = 248 & 490;
  assign n357 = 316 & n356;
  assign n358 = 251 & 490;
  assign n359 = ~316 & n358;
  assign n360 = ~n357 & ~n359;
  assign n361 = 242 & 316;
  assign n362 = 254 & ~316;
  assign n363 = ~n361 & ~n362;
  assign n364 = ~490 & n363;
  assign n365 = n360 & ~n364;
  assign n366 = 248 & 479;
  assign n367 = 308 & n366;
  assign n368 = 251 & 479;
  assign n369 = ~308 & n368;
  assign n370 = ~n367 & ~n369;
  assign n371 = 242 & 308;
  assign n372 = 254 & ~308;
  assign n373 = ~n371 & ~n372;
  assign n374 = ~479 & n373;
  assign n375 = n370 & ~n374;
  assign n376 = 248 & 302;
  assign n377 = 251 & ~302;
  assign n378 = ~n376 & ~n377;
  assign n379 = 242 & 293;
  assign n380 = 254 & ~293;
  assign n381 = ~n379 & ~n380;
  assign n382 = ~n365 & ~n375;
  assign n383 = ~n378 & n382;
  assign n384 = n381 & n383;
  assign n385 = 534 & ~598;
  assign n386 = 351 & n385;
  assign n387 = 534 & ~597;
  assign n388 = ~351 & n387;
  assign n389 = ~n386 & ~n388;
  assign n390 = 351 & ~595;
  assign n391 = ~351 & ~596;
  assign n392 = ~n390 & ~n391;
  assign n393 = ~534 & n392;
  assign n394 = n389 & ~n393;
  assign n395 = 523 & ~598;
  assign n396 = 341 & n395;
  assign n397 = 523 & ~597;
  assign n398 = ~341 & n397;
  assign n399 = ~n396 & ~n398;
  assign n400 = 341 & ~595;
  assign n401 = ~341 & ~596;
  assign n402 = ~n400 & ~n401;
  assign n403 = ~523 & n402;
  assign n404 = n399 & ~n403;
  assign n405 = 514 & ~598;
  assign n406 = ~514 & 595;
  assign n407 = ~n405 & ~n406;
  assign n408 = 503 & ~598;
  assign n409 = 324 & n408;
  assign n410 = 503 & ~597;
  assign n411 = ~324 & n410;
  assign n412 = ~n409 & ~n411;
  assign n413 = 324 & ~595;
  assign n414 = ~324 & ~596;
  assign n415 = ~n413 & ~n414;
  assign n416 = ~503 & n415;
  assign n417 = n412 & ~n416;
  assign n418 = ~n394 & ~n404;
  assign n419 = ~n407 & n418;
  assign n420 = ~n417 & n419;
  assign n421 = 248 & 361;
  assign n422 = 251 & ~361;
  assign n423 = ~n421 & ~n422;
  assign n424 = n384 & n420;
  assign 5240 = ~n423 & n424;
  assign n426 = 435 & ~598;
  assign n427 = 234 & n426;
  assign n428 = 435 & ~597;
  assign n429 = ~234 & n428;
  assign n430 = ~n427 & ~n429;
  assign n431 = 234 & ~595;
  assign n432 = ~234 & ~596;
  assign n433 = ~n431 & ~n432;
  assign n434 = ~435 & n433;
  assign n435 = n430 & ~n434;
  assign n436 = 422 & ~598;
  assign n437 = 226 & n436;
  assign n438 = 422 & ~597;
  assign n439 = ~226 & n438;
  assign n440 = ~n437 & ~n439;
  assign n441 = 226 & ~595;
  assign n442 = ~226 & ~596;
  assign n443 = ~n441 & ~n442;
  assign n444 = ~422 & n443;
  assign n445 = n440 & ~n444;
  assign n446 = 468 & ~598;
  assign n447 = 218 & n446;
  assign n448 = 468 & ~597;
  assign n449 = ~218 & n448;
  assign n450 = ~n447 & ~n449;
  assign n451 = 218 & ~595;
  assign n452 = ~218 & ~596;
  assign n453 = ~n451 & ~n452;
  assign n454 = ~468 & n453;
  assign n455 = n450 & ~n454;
  assign n456 = 457 & ~598;
  assign n457 = 210 & n456;
  assign n458 = 457 & ~597;
  assign n459 = ~210 & n458;
  assign n460 = ~n457 & ~n459;
  assign n461 = 210 & ~595;
  assign n462 = ~210 & ~596;
  assign n463 = ~n461 & ~n462;
  assign n464 = ~457 & n463;
  assign n465 = n460 & ~n464;
  assign n466 = ~n435 & ~n445;
  assign n467 = ~n455 & n466;
  assign n468 = ~n465 & n467;
  assign n469 = 374 & ~598;
  assign n470 = 281 & n469;
  assign n471 = 374 & ~597;
  assign n472 = ~281 & n471;
  assign n473 = ~n470 & ~n472;
  assign n474 = 281 & ~595;
  assign n475 = ~281 & ~596;
  assign n476 = ~n474 & ~n475;
  assign n477 = ~374 & n476;
  assign n478 = n473 & ~n477;
  assign n479 = 411 & ~598;
  assign n480 = 273 & n479;
  assign n481 = 411 & ~597;
  assign n482 = ~273 & n481;
  assign n483 = ~n480 & ~n482;
  assign n484 = 273 & ~595;
  assign n485 = ~273 & ~596;
  assign n486 = ~n484 & ~n485;
  assign n487 = ~411 & n486;
  assign n488 = n483 & ~n487;
  assign n489 = 400 & ~598;
  assign n490 = 265 & n489;
  assign n491 = 400 & ~597;
  assign n492 = ~265 & n491;
  assign n493 = ~n490 & ~n492;
  assign n494 = 265 & ~595;
  assign n495 = ~265 & ~596;
  assign n496 = ~n494 & ~n495;
  assign n497 = ~400 & n496;
  assign n498 = n493 & ~n497;
  assign n499 = 389 & ~598;
  assign n500 = 257 & n499;
  assign n501 = 389 & ~597;
  assign n502 = ~257 & n501;
  assign n503 = ~n500 & ~n502;
  assign n504 = 257 & ~595;
  assign n505 = ~257 & ~596;
  assign n506 = ~n504 & ~n505;
  assign n507 = ~389 & n506;
  assign n508 = n503 & ~n507;
  assign n509 = ~n478 & ~n488;
  assign n510 = ~n498 & n509;
  assign n511 = ~n508 & n510;
  assign n512 = 248 & 446;
  assign n513 = 206 & n512;
  assign n514 = 251 & 446;
  assign n515 = ~206 & n514;
  assign n516 = ~n513 & ~n515;
  assign n517 = 206 & 242;
  assign n518 = ~206 & 254;
  assign n519 = ~n517 & ~n518;
  assign n520 = ~446 & n519;
  assign n521 = n516 & ~n520;
  assign n522 = n468 & n511;
  assign 5388 = ~n521 & n522;
  assign n524 = 226 & ~335;
  assign n525 = 233 & 335;
  assign n526 = ~n524 & ~n525;
  assign n527 = ~422 & ~n526;
  assign n528 = 422 & n526;
  assign n529 = ~n527 & ~n528;
  assign n530 = 218 & ~335;
  assign n531 = 225 & 335;
  assign n532 = ~n530 & ~n531;
  assign n533 = ~468 & ~n532;
  assign n534 = 468 & n532;
  assign n535 = ~n533 & ~n534;
  assign n536 = 210 & ~335;
  assign n537 = 217 & 335;
  assign n538 = ~n536 & ~n537;
  assign n539 = ~457 & ~n538;
  assign n540 = 457 & n538;
  assign n541 = ~n539 & ~n540;
  assign n542 = 206 & ~335;
  assign n543 = 209 & 335;
  assign n544 = ~n542 & ~n543;
  assign n545 = ~446 & ~n544;
  assign n546 = 446 & n544;
  assign n547 = ~n545 & ~n546;
  assign n548 = ~n529 & ~n535;
  assign n549 = ~n541 & n548;
  assign n550 = ~n547 & n549;
  assign n551 = 281 & ~335;
  assign n552 = 288 & 335;
  assign n553 = ~n551 & ~n552;
  assign n554 = ~374 & ~n553;
  assign n555 = 374 & n553;
  assign n556 = ~n554 & ~n555;
  assign n557 = 273 & ~335;
  assign n558 = 280 & 335;
  assign n559 = ~n557 & ~n558;
  assign n560 = ~411 & ~n559;
  assign n561 = 411 & n559;
  assign n562 = ~n560 & ~n561;
  assign n563 = 265 & ~335;
  assign n564 = 272 & 335;
  assign n565 = ~n563 & ~n564;
  assign n566 = ~400 & ~n565;
  assign n567 = 400 & n565;
  assign n568 = ~n566 & ~n567;
  assign n569 = 257 & ~335;
  assign n570 = 264 & 335;
  assign n571 = ~n569 & ~n570;
  assign n572 = ~389 & ~n571;
  assign n573 = 389 & n571;
  assign n574 = ~n572 & ~n573;
  assign n575 = 234 & ~335;
  assign n576 = 241 & 335;
  assign n577 = ~n575 & ~n576;
  assign n578 = ~435 & ~n577;
  assign n579 = 435 & n577;
  assign n580 = ~n578 & ~n579;
  assign n581 = ~n556 & ~n562;
  assign n582 = ~n568 & n581;
  assign n583 = ~n574 & n582;
  assign n584 = ~n580 & n583;
  assign 6641 = n550 & n584;
  assign n586 = 302 & ~332;
  assign n587 = 307 & 332;
  assign n588 = ~n586 & ~n587;
  assign n589 = 316 & ~332;
  assign n590 = 323 & 332;
  assign n591 = ~n589 & ~n590;
  assign n592 = 490 & n591;
  assign n593 = ~490 & ~n591;
  assign n594 = ~n592 & ~n593;
  assign n595 = 308 & ~332;
  assign n596 = 315 & 332;
  assign n597 = ~n595 & ~n596;
  assign n598 = 479 & n597;
  assign n599 = ~479 & ~n597;
  assign n600 = ~n598 & ~n599;
  assign n601 = 293 & ~332;
  assign n602 = 299 & 332;
  assign n603 = ~n601 & ~n602;
  assign n604 = n588 & ~n594;
  assign n605 = ~n600 & n604;
  assign n606 = n603 & n605;
  assign n607 = 332 & 338;
  assign n608 = 332 & ~n607;
  assign n609 = 514 & n608;
  assign n610 = ~514 & ~n608;
  assign n611 = ~n609 & ~n610;
  assign n612 = ~332 & 361;
  assign n613 = 332 & 366;
  assign n614 = ~n612 & ~n613;
  assign n615 = ~332 & 341;
  assign n616 = 332 & 348;
  assign n617 = ~n615 & ~n616;
  assign n618 = 523 & n617;
  assign n619 = ~523 & ~n617;
  assign n620 = ~n618 & ~n619;
  assign n621 = 324 & ~332;
  assign n622 = 331 & 332;
  assign n623 = ~n621 & ~n622;
  assign n624 = 503 & n623;
  assign n625 = ~503 & ~n623;
  assign n626 = ~n624 & ~n625;
  assign n627 = ~332 & 351;
  assign n628 = 332 & 358;
  assign n629 = ~n627 & ~n628;
  assign n630 = 534 & n629;
  assign n631 = ~534 & ~n629;
  assign n632 = ~n630 & ~n631;
  assign n633 = ~n611 & n614;
  assign n634 = ~n620 & n633;
  assign n635 = ~n626 & n634;
  assign n636 = ~n632 & n635;
  assign 6643 = n606 & n636;
  assign n638 = ~n594 & ~n600;
  assign n639 = n588 & n638;
  assign n640 = n603 & n639;
  assign n641 = n614 & ~n632;
  assign n642 = ~n620 & n641;
  assign n643 = ~n611 & n642;
  assign n644 = ~n626 & n643;
  assign 6646 = n640 & n644;
  assign n646 = ~n529 & ~n541;
  assign n647 = ~n535 & n646;
  assign n648 = ~n547 & n647;
  assign n649 = ~n556 & ~n574;
  assign n650 = ~n568 & n649;
  assign n651 = ~n580 & n650;
  assign n652 = ~n562 & n651;
  assign 6648 = n648 & n652;
  assign n654 = ~308 & 316;
  assign n655 = 308 & ~316;
  assign n656 = ~n654 & ~n655;
  assign n657 = ~293 & 302;
  assign n658 = 293 & ~302;
  assign n659 = ~n657 & ~n658;
  assign n660 = ~n656 & n659;
  assign n661 = n656 & ~n659;
  assign n662 = ~n660 & ~n661;
  assign n663 = ~361 & 369;
  assign n664 = 361 & ~369;
  assign n665 = ~n663 & ~n664;
  assign n666 = ~341 & 351;
  assign n667 = 341 & ~351;
  assign n668 = ~n666 & ~n667;
  assign n669 = ~n665 & n668;
  assign n670 = 324 & n669;
  assign n671 = n665 & n668;
  assign n672 = ~324 & n671;
  assign n673 = ~n670 & ~n672;
  assign n674 = n665 & ~n668;
  assign n675 = 324 & n674;
  assign n676 = ~n665 & ~n668;
  assign n677 = ~324 & n676;
  assign n678 = ~n675 & ~n677;
  assign n679 = n673 & n678;
  assign n680 = ~n662 & n679;
  assign n681 = n662 & ~n679;
  assign 6716 = n680 | n681;
  assign n683 = ~218 & 226;
  assign n684 = 218 & ~226;
  assign n685 = ~n683 & ~n684;
  assign n686 = ~206 & 210;
  assign n687 = 206 & ~210;
  assign n688 = ~n686 & ~n687;
  assign n689 = ~n685 & n688;
  assign n690 = n685 & ~n688;
  assign n691 = ~n689 & ~n690;
  assign n692 = ~281 & 289;
  assign n693 = 281 & ~289;
  assign n694 = ~n692 & ~n693;
  assign n695 = ~265 & 273;
  assign n696 = 265 & ~273;
  assign n697 = ~n695 & ~n696;
  assign n698 = ~234 & 257;
  assign n699 = 234 & ~257;
  assign n700 = ~n698 & ~n699;
  assign n701 = ~n694 & n697;
  assign n702 = n700 & n701;
  assign n703 = n694 & n697;
  assign n704 = ~n700 & n703;
  assign n705 = ~n702 & ~n704;
  assign n706 = n694 & ~n697;
  assign n707 = n700 & n706;
  assign n708 = ~n694 & ~n697;
  assign n709 = ~n700 & n708;
  assign n710 = ~n707 & ~n709;
  assign n711 = n705 & n710;
  assign n712 = ~n691 & n711;
  assign n713 = n691 & ~n711;
  assign 6877 = n712 | n713;
  assign n715 = 446 & ~n544;
  assign n716 = 457 & ~n538;
  assign n717 = ~n547 & n716;
  assign n718 = 468 & ~n532;
  assign n719 = ~n541 & ~n547;
  assign n720 = n718 & n719;
  assign n721 = 422 & ~n526;
  assign n722 = ~n535 & ~n547;
  assign n723 = n721 & n722;
  assign n724 = ~n541 & n723;
  assign n725 = ~n715 & ~n717;
  assign n726 = ~n720 & n725;
  assign n727 = ~n724 & n726;
  assign n728 = 435 & ~n577;
  assign n729 = 389 & ~n571;
  assign n730 = ~n580 & n729;
  assign n731 = 400 & ~n565;
  assign n732 = ~n574 & ~n580;
  assign n733 = n731 & n732;
  assign n734 = 411 & ~n559;
  assign n735 = ~n568 & ~n580;
  assign n736 = n734 & n735;
  assign n737 = ~n574 & n736;
  assign n738 = 374 & ~n553;
  assign n739 = ~n562 & ~n568;
  assign n740 = ~n580 & n739;
  assign n741 = n738 & n740;
  assign n742 = ~n574 & n741;
  assign n743 = ~n728 & ~n730;
  assign n744 = ~n733 & n743;
  assign n745 = ~n737 & n744;
  assign n746 = ~n742 & n745;
  assign n747 = n550 & ~n746;
  assign 6924 = ~n727 | n747;
  assign n749 = ~n588 & n603;
  assign n750 = 479 & ~n597;
  assign n751 = n588 & n603;
  assign n752 = n750 & n751;
  assign n753 = 490 & ~n591;
  assign n754 = ~n600 & n603;
  assign n755 = n753 & n754;
  assign n756 = n588 & n755;
  assign n757 = n603 & ~n749;
  assign n758 = ~n752 & n757;
  assign n759 = ~n756 & n758;
  assign n760 = 503 & ~n623;
  assign n761 = 514 & ~n608;
  assign n762 = ~n626 & n761;
  assign n763 = 523 & ~n617;
  assign n764 = ~n611 & ~n626;
  assign n765 = n763 & n764;
  assign n766 = 534 & ~n629;
  assign n767 = ~n620 & ~n626;
  assign n768 = n766 & n767;
  assign n769 = ~n611 & n768;
  assign n770 = ~n620 & ~n632;
  assign n771 = ~n626 & n770;
  assign n772 = ~n614 & n771;
  assign n773 = ~n611 & n772;
  assign n774 = ~n760 & ~n762;
  assign n775 = ~n765 & n774;
  assign n776 = ~n769 & n775;
  assign n777 = ~n773 & n776;
  assign n778 = n606 & ~n777;
  assign 6925 = ~n759 | n778;
  assign n780 = n648 & ~n746;
  assign 6926 = ~n727 | n780;
  assign n782 = n640 & ~n777;
  assign 6927 = ~n759 | n782;
  assign n784 = ~619 & n423;
  assign n785 = ~625 & n784;
  assign n786 = ~54 & n614;
  assign n787 = 54 & ~n614;
  assign n788 = ~n786 & ~n787;
  assign n789 = 619 & ~n788;
  assign n790 = ~625 & n789;
  assign n791 = 131 & ~619;
  assign n792 = 625 & n791;
  assign n793 = ~n785 & ~n790;
  assign 7015 = ~n792 & n793;
  assign n795 = ~619 & n394;
  assign n796 = ~625 & n795;
  assign n797 = 54 & n614;
  assign n798 = n614 & ~n797;
  assign n799 = ~n632 & n798;
  assign n800 = n632 & ~n798;
  assign n801 = ~n799 & ~n800;
  assign n802 = 619 & ~n801;
  assign n803 = ~625 & n802;
  assign n804 = 129 & ~619;
  assign n805 = 625 & n804;
  assign n806 = ~n796 & ~n803;
  assign 7363 = ~n805 & n806;
  assign n808 = ~619 & n478;
  assign n809 = ~625 & n808;
  assign n810 = ~4 & ~n556;
  assign n811 = 4 & n556;
  assign n812 = ~n810 & ~n811;
  assign n813 = 619 & ~n812;
  assign n814 = ~625 & n813;
  assign n815 = 117 & ~619;
  assign n816 = 625 & n815;
  assign n817 = ~n809 & ~n814;
  assign 7365 = ~n816 & n817;
  assign n819 = n588 & n750;
  assign n820 = ~n600 & n753;
  assign n821 = n588 & n820;
  assign n822 = n588 & ~n819;
  assign n823 = ~n821 & n822;
  assign n824 = n603 & ~n823;
  assign n825 = ~n603 & n823;
  assign n826 = ~n824 & ~n825;
  assign n827 = 54 & n636;
  assign n828 = n777 & ~n827;
  assign n829 = n826 & n828;
  assign n830 = ~n639 & n823;
  assign n831 = n603 & n830;
  assign n832 = ~n603 & ~n830;
  assign n833 = ~n831 & ~n832;
  assign n834 = ~n828 & ~n833;
  assign 7432 = ~n829 & ~n834;
  assign n836 = ~610 & ~7015;
  assign n837 = ~607 & n836;
  assign n838 = 610 & ~7365;
  assign n839 = ~607 & n838;
  assign n840 = 11 & ~610;
  assign n841 = 607 & n840;
  assign n842 = 61 & 610;
  assign n843 = 607 & n842;
  assign n844 = ~n837 & ~n839;
  assign n845 = ~n841 & n844;
  assign 7449 = n843 | ~n845;
  assign n847 = ~619 & n417;
  assign n848 = ~625 & n847;
  assign n849 = ~n611 & n763;
  assign n850 = ~n620 & n766;
  assign n851 = ~n611 & n850;
  assign n852 = ~n614 & n770;
  assign n853 = ~n611 & n852;
  assign n854 = ~n620 & n797;
  assign n855 = ~n632 & n854;
  assign n856 = ~n611 & n855;
  assign n857 = ~n761 & ~n849;
  assign n858 = ~n851 & n857;
  assign n859 = ~n853 & n858;
  assign n860 = ~n856 & n859;
  assign n861 = ~n626 & n860;
  assign n862 = n626 & ~n860;
  assign n863 = ~n861 & ~n862;
  assign n864 = 619 & ~n863;
  assign n865 = ~625 & n864;
  assign n866 = 52 & ~619;
  assign n867 = 625 & n866;
  assign n868 = ~n848 & ~n865;
  assign 7465 = ~n867 & n868;
  assign n870 = ~619 & n407;
  assign n871 = ~625 & n870;
  assign n872 = ~n763 & ~n850;
  assign n873 = ~n852 & n872;
  assign n874 = ~n855 & n873;
  assign n875 = ~n611 & n874;
  assign n876 = n611 & ~n874;
  assign n877 = ~n875 & ~n876;
  assign n878 = 619 & ~n877;
  assign n879 = ~625 & n878;
  assign n880 = 130 & ~619;
  assign n881 = 625 & n880;
  assign n882 = ~n871 & ~n879;
  assign 7466 = ~n881 & n882;
  assign n884 = ~619 & n404;
  assign n885 = ~625 & n884;
  assign n886 = ~n614 & ~n632;
  assign n887 = ~n632 & n797;
  assign n888 = ~n766 & ~n886;
  assign n889 = ~n887 & n888;
  assign n890 = ~n620 & n889;
  assign n891 = n620 & ~n889;
  assign n892 = ~n890 & ~n891;
  assign n893 = 619 & ~n892;
  assign n894 = ~625 & n893;
  assign n895 = 119 & ~619;
  assign n896 = 625 & n895;
  assign n897 = ~n885 & ~n894;
  assign 7467 = ~n896 & n897;
  assign n899 = ~613 & ~7015;
  assign n900 = ~616 & n899;
  assign n901 = 613 & ~7365;
  assign n902 = ~616 & n901;
  assign n903 = 11 & ~613;
  assign n904 = 616 & n903;
  assign n905 = 61 & 613;
  assign n906 = 616 & n905;
  assign n907 = ~n900 & ~n902;
  assign n908 = ~n904 & n907;
  assign 7469 = n906 | ~n908;
  assign n910 = ~619 & n435;
  assign n911 = ~625 & n910;
  assign n912 = ~n574 & n731;
  assign n913 = ~n568 & n734;
  assign n914 = ~n574 & n913;
  assign n915 = n738 & n739;
  assign n916 = ~n574 & n915;
  assign n917 = 4 & ~n556;
  assign n918 = ~n568 & n917;
  assign n919 = ~n562 & n918;
  assign n920 = ~n574 & n919;
  assign n921 = ~n729 & ~n912;
  assign n922 = ~n914 & n921;
  assign n923 = ~n916 & n922;
  assign n924 = ~n920 & n923;
  assign n925 = ~n580 & n924;
  assign n926 = n580 & ~n924;
  assign n927 = ~n925 & ~n926;
  assign n928 = 619 & ~n927;
  assign n929 = ~625 & n928;
  assign n930 = 122 & ~619;
  assign n931 = 625 & n930;
  assign n932 = ~n911 & ~n929;
  assign 7470 = ~n931 & n932;
  assign n934 = ~619 & n508;
  assign n935 = ~625 & n934;
  assign n936 = ~n731 & ~n913;
  assign n937 = ~n915 & n936;
  assign n938 = ~n919 & n937;
  assign n939 = ~n574 & n938;
  assign n940 = n574 & ~n938;
  assign n941 = ~n939 & ~n940;
  assign n942 = 619 & ~n941;
  assign n943 = ~625 & n942;
  assign n944 = 128 & ~619;
  assign n945 = 625 & n944;
  assign n946 = ~n935 & ~n943;
  assign 7471 = ~n945 & n946;
  assign n948 = ~619 & n498;
  assign n949 = ~625 & n948;
  assign n950 = ~n562 & n738;
  assign n951 = ~n562 & n917;
  assign n952 = ~n734 & ~n950;
  assign n953 = ~n951 & n952;
  assign n954 = ~n568 & n953;
  assign n955 = n568 & ~n953;
  assign n956 = ~n954 & ~n955;
  assign n957 = 619 & ~n956;
  assign n958 = ~625 & n957;
  assign n959 = 127 & ~619;
  assign n960 = 625 & n959;
  assign n961 = ~n949 & ~n958;
  assign 7472 = ~n960 & n961;
  assign n963 = ~619 & n488;
  assign n964 = ~625 & n963;
  assign n965 = ~n738 & ~n917;
  assign n966 = ~n562 & n965;
  assign n967 = n562 & ~n965;
  assign n968 = ~n966 & ~n967;
  assign n969 = 619 & ~n968;
  assign n970 = ~625 & n969;
  assign n971 = 126 & ~619;
  assign n972 = 625 & n971;
  assign n973 = ~n964 & ~n970;
  assign 7473 = ~n972 & n973;
  assign n975 = ~n591 & n597;
  assign n976 = n591 & ~n597;
  assign n977 = ~n975 & ~n976;
  assign n978 = n588 & ~n603;
  assign n979 = ~n749 & ~n978;
  assign n980 = ~n977 & n979;
  assign n981 = n977 & ~n979;
  assign n982 = ~n980 & ~n981;
  assign n983 = ~n617 & n629;
  assign n984 = n617 & ~n629;
  assign n985 = ~n983 & ~n984;
  assign n986 = ~332 & 369;
  assign n987 = 332 & 372;
  assign n988 = ~n986 & ~n987;
  assign n989 = ~n614 & n988;
  assign n990 = n614 & ~n988;
  assign n991 = ~n989 & ~n990;
  assign n992 = ~n608 & n623;
  assign n993 = n608 & ~n623;
  assign n994 = ~n992 & ~n993;
  assign n995 = ~n985 & n991;
  assign n996 = n994 & n995;
  assign n997 = n985 & n991;
  assign n998 = ~n994 & n997;
  assign n999 = ~n996 & ~n998;
  assign n1000 = n985 & ~n991;
  assign n1001 = n994 & n1000;
  assign n1002 = ~n985 & ~n991;
  assign n1003 = ~n994 & n1002;
  assign n1004 = ~n1001 & ~n1003;
  assign n1005 = n999 & n1004;
  assign n1006 = ~n982 & n1005;
  assign n1007 = n982 & ~n1005;
  assign 7474 = n1006 | n1007;
  assign n1009 = ~n553 & n559;
  assign n1010 = n553 & ~n559;
  assign n1011 = ~n1009 & ~n1010;
  assign n1012 = ~n565 & n571;
  assign n1013 = n565 & ~n571;
  assign n1014 = ~n1012 & ~n1013;
  assign n1015 = ~n1011 & n1014;
  assign n1016 = n1011 & ~n1014;
  assign n1017 = ~n1015 & ~n1016;
  assign n1018 = n526 & ~n577;
  assign n1019 = ~n526 & n577;
  assign n1020 = ~n1018 & ~n1019;
  assign n1021 = ~n532 & n538;
  assign n1022 = n532 & ~n538;
  assign n1023 = ~n1021 & ~n1022;
  assign n1024 = 289 & ~335;
  assign n1025 = 292 & 335;
  assign n1026 = ~n1024 & ~n1025;
  assign n1027 = ~n544 & n1026;
  assign n1028 = n544 & ~n1026;
  assign n1029 = ~n1027 & ~n1028;
  assign n1030 = ~n1020 & n1023;
  assign n1031 = n1029 & n1030;
  assign n1032 = n1020 & n1023;
  assign n1033 = ~n1029 & n1032;
  assign n1034 = ~n1031 & ~n1033;
  assign n1035 = n1020 & ~n1023;
  assign n1036 = n1029 & n1035;
  assign n1037 = ~n1020 & ~n1023;
  assign n1038 = ~n1029 & n1037;
  assign n1039 = ~n1036 & ~n1038;
  assign n1040 = n1034 & n1039;
  assign n1041 = ~n1017 & n1040;
  assign n1042 = n1017 & ~n1040;
  assign 7476 = n1041 | n1042;
  assign n1044 = 4 & n652;
  assign n1045 = n746 & ~n1044;
  assign n1046 = ~n529 & n1045;
  assign n1047 = n529 & ~n1045;
  assign n1048 = ~n1046 & ~n1047;
  assign n1049 = ~n535 & ~n721;
  assign n1050 = n535 & n721;
  assign n1051 = ~n1049 & ~n1050;
  assign n1052 = n1045 & ~n1051;
  assign n1053 = ~422 & n526;
  assign n1054 = ~n535 & ~n1053;
  assign n1055 = n535 & n1053;
  assign n1056 = ~n1054 & ~n1055;
  assign n1057 = ~n1045 & n1056;
  assign n1058 = ~n1052 & ~n1057;
  assign n1059 = ~n535 & n721;
  assign n1060 = ~n718 & ~n1059;
  assign n1061 = ~n541 & ~n1060;
  assign n1062 = n541 & n1060;
  assign n1063 = ~n1061 & ~n1062;
  assign n1064 = n1045 & n1063;
  assign n1065 = ~n548 & n1060;
  assign n1066 = ~n541 & n1065;
  assign n1067 = n541 & ~n1065;
  assign n1068 = ~n1066 & ~n1067;
  assign n1069 = ~n1045 & ~n1068;
  assign n1070 = ~n1064 & ~n1069;
  assign n1071 = ~n541 & n718;
  assign n1072 = ~n541 & n1059;
  assign n1073 = ~n716 & ~n1071;
  assign n1074 = ~n1072 & n1073;
  assign n1075 = ~n547 & ~n1074;
  assign n1076 = n547 & n1074;
  assign n1077 = ~n1075 & ~n1076;
  assign n1078 = n1045 & n1077;
  assign n1079 = ~n549 & n1074;
  assign n1080 = ~n547 & n1079;
  assign n1081 = n547 & ~n1079;
  assign n1082 = ~n1080 & ~n1081;
  assign n1083 = ~n1045 & ~n1082;
  assign n1084 = ~n1078 & ~n1083;
  assign n1085 = n812 & n968;
  assign n1086 = n956 & n1085;
  assign n1087 = n941 & n1086;
  assign n1088 = n927 & n1087;
  assign n1089 = n1048 & n1088;
  assign n1090 = n1058 & n1089;
  assign n1091 = n1070 & n1090;
  assign 7503 = n1084 & n1091;
  assign n1093 = ~n594 & n828;
  assign n1094 = n594 & ~n828;
  assign n1095 = ~n1093 & ~n1094;
  assign n1096 = ~n600 & ~n753;
  assign n1097 = n600 & n753;
  assign n1098 = ~n1096 & ~n1097;
  assign n1099 = n828 & ~n1098;
  assign n1100 = ~490 & n591;
  assign n1101 = ~n600 & ~n1100;
  assign n1102 = n600 & n1100;
  assign n1103 = ~n1101 & ~n1102;
  assign n1104 = ~n828 & n1103;
  assign n1105 = ~n1099 & ~n1104;
  assign n1106 = ~n750 & ~n820;
  assign n1107 = n588 & ~n1106;
  assign n1108 = ~n588 & n1106;
  assign n1109 = ~n1107 & ~n1108;
  assign n1110 = n828 & n1109;
  assign n1111 = ~n638 & n1106;
  assign n1112 = n588 & n1111;
  assign n1113 = ~n588 & ~n1111;
  assign n1114 = ~n1112 & ~n1113;
  assign n1115 = ~n828 & ~n1114;
  assign n1116 = ~n1110 & ~n1115;
  assign n1117 = n788 & n801;
  assign n1118 = n892 & n1117;
  assign n1119 = n877 & n1118;
  assign n1120 = n863 & n1119;
  assign n1121 = n1095 & n1120;
  assign n1122 = n1105 & n1121;
  assign n1123 = n1116 & n1122;
  assign 7504 = 7432 & n1123;
  assign n1125 = ~571 & ~7015;
  assign n1126 = ~574 & n1125;
  assign n1127 = 571 & ~7365;
  assign n1128 = ~574 & n1127;
  assign n1129 = 182 & ~571;
  assign n1130 = 574 & n1129;
  assign n1131 = 185 & 571;
  assign n1132 = 574 & n1131;
  assign n1133 = ~n1126 & ~n1128;
  assign n1134 = ~n1130 & n1133;
  assign n1135 = ~n1132 & n1134;
  assign 7506 = 137 & ~n1135;
  assign n1137 = ~577 & ~7015;
  assign n1138 = ~580 & n1137;
  assign n1139 = 577 & ~7365;
  assign n1140 = ~580 & n1139;
  assign n1141 = 182 & ~577;
  assign n1142 = 580 & n1141;
  assign n1143 = 185 & 577;
  assign n1144 = 580 & n1143;
  assign n1145 = ~n1138 & ~n1140;
  assign n1146 = ~n1142 & n1145;
  assign n1147 = ~n1144 & n1146;
  assign 7511 = 137 & ~n1147;
  assign n1149 = ~610 & ~7465;
  assign n1150 = ~607 & n1149;
  assign n1151 = 610 & ~7470;
  assign n1152 = ~607 & n1151;
  assign n1153 = 43 & ~610;
  assign n1154 = 607 & n1153;
  assign n1155 = 37 & 610;
  assign n1156 = 607 & n1155;
  assign n1157 = ~n1150 & ~n1152;
  assign n1158 = ~n1154 & n1157;
  assign 7515 = n1156 | ~n1158;
  assign n1160 = ~610 & ~7466;
  assign n1161 = ~607 & n1160;
  assign n1162 = 610 & ~7471;
  assign n1163 = ~607 & n1162;
  assign n1164 = 76 & ~610;
  assign n1165 = 607 & n1164;
  assign n1166 = 20 & 610;
  assign n1167 = 607 & n1166;
  assign n1168 = ~n1161 & ~n1163;
  assign n1169 = ~n1165 & n1168;
  assign 7516 = n1167 | ~n1169;
  assign n1171 = ~610 & ~7467;
  assign n1172 = ~607 & n1171;
  assign n1173 = 610 & ~7472;
  assign n1174 = ~607 & n1173;
  assign n1175 = 73 & ~610;
  assign n1176 = 607 & n1175;
  assign n1177 = 17 & 610;
  assign n1178 = 607 & n1177;
  assign n1179 = ~n1172 & ~n1174;
  assign n1180 = ~n1176 & n1179;
  assign 7517 = n1178 | ~n1180;
  assign n1182 = ~610 & ~7363;
  assign n1183 = ~607 & n1182;
  assign n1184 = 610 & ~7473;
  assign n1185 = ~607 & n1184;
  assign n1186 = 67 & ~610;
  assign n1187 = 607 & n1186;
  assign n1188 = 70 & 610;
  assign n1189 = 607 & n1188;
  assign n1190 = ~n1183 & ~n1185;
  assign n1191 = ~n1187 & n1190;
  assign 7518 = n1189 | ~n1191;
  assign n1193 = ~613 & ~7465;
  assign n1194 = ~616 & n1193;
  assign n1195 = 613 & ~7470;
  assign n1196 = ~616 & n1195;
  assign n1197 = 43 & ~613;
  assign n1198 = 616 & n1197;
  assign n1199 = 37 & 613;
  assign n1200 = 616 & n1199;
  assign n1201 = ~n1194 & ~n1196;
  assign n1202 = ~n1198 & n1201;
  assign 7519 = n1200 | ~n1202;
  assign n1204 = ~613 & ~7466;
  assign n1205 = ~616 & n1204;
  assign n1206 = 613 & ~7471;
  assign n1207 = ~616 & n1206;
  assign n1208 = 76 & ~613;
  assign n1209 = 616 & n1208;
  assign n1210 = 20 & 613;
  assign n1211 = 616 & n1210;
  assign n1212 = ~n1205 & ~n1207;
  assign n1213 = ~n1209 & n1212;
  assign 7520 = n1211 | ~n1213;
  assign n1215 = ~613 & ~7467;
  assign n1216 = ~616 & n1215;
  assign n1217 = 613 & ~7472;
  assign n1218 = ~616 & n1217;
  assign n1219 = 73 & ~613;
  assign n1220 = 616 & n1219;
  assign n1221 = 17 & 613;
  assign n1222 = 616 & n1221;
  assign n1223 = ~n1216 & ~n1218;
  assign n1224 = ~n1220 & n1223;
  assign 7521 = n1222 | ~n1224;
  assign n1226 = ~613 & ~7363;
  assign n1227 = ~616 & n1226;
  assign n1228 = 613 & ~7473;
  assign n1229 = ~616 & n1228;
  assign n1230 = 67 & ~613;
  assign n1231 = 616 & n1230;
  assign n1232 = 70 & 613;
  assign n1233 = 616 & n1232;
  assign n1234 = ~n1227 & ~n1229;
  assign n1235 = ~n1231 & n1234;
  assign 7522 = n1233 | ~n1235;
  assign n1237 = ~571 & ~7465;
  assign n1238 = ~574 & n1237;
  assign n1239 = 571 & ~7470;
  assign n1240 = ~574 & n1239;
  assign n1241 = 200 & ~571;
  assign n1242 = 574 & n1241;
  assign n1243 = 170 & 571;
  assign n1244 = 574 & n1243;
  assign n1245 = ~n1238 & ~n1240;
  assign n1246 = ~n1242 & n1245;
  assign n1247 = ~n1244 & n1246;
  assign 7600 = 137 & ~n1247;
  assign n1249 = ~571 & ~7363;
  assign n1250 = ~574 & n1249;
  assign n1251 = 571 & ~7473;
  assign n1252 = ~574 & n1251;
  assign n1253 = 188 & ~571;
  assign n1254 = 574 & n1253;
  assign n1255 = 158 & 571;
  assign n1256 = 574 & n1255;
  assign n1257 = ~n1250 & ~n1252;
  assign n1258 = ~n1254 & n1257;
  assign n1259 = ~n1256 & n1258;
  assign 7601 = 137 & ~n1259;
  assign n1261 = ~571 & ~7467;
  assign n1262 = ~574 & n1261;
  assign n1263 = 571 & ~7472;
  assign n1264 = ~574 & n1263;
  assign n1265 = 155 & ~571;
  assign n1266 = 574 & n1265;
  assign n1267 = 152 & 571;
  assign n1268 = 574 & n1267;
  assign n1269 = ~n1262 & ~n1264;
  assign n1270 = ~n1266 & n1269;
  assign n1271 = ~n1268 & n1270;
  assign 7602 = 137 & ~n1271;
  assign n1273 = ~571 & ~7466;
  assign n1274 = ~574 & n1273;
  assign n1275 = 571 & ~7471;
  assign n1276 = ~574 & n1275;
  assign n1277 = 149 & ~571;
  assign n1278 = 574 & n1277;
  assign n1279 = 146 & 571;
  assign n1280 = 574 & n1279;
  assign n1281 = ~n1274 & ~n1276;
  assign n1282 = ~n1278 & n1281;
  assign n1283 = ~n1280 & n1282;
  assign 7603 = 137 & ~n1283;
  assign n1285 = ~577 & ~7465;
  assign n1286 = ~580 & n1285;
  assign n1287 = 577 & ~7470;
  assign n1288 = ~580 & n1287;
  assign n1289 = 200 & ~577;
  assign n1290 = 580 & n1289;
  assign n1291 = 170 & 577;
  assign n1292 = 580 & n1291;
  assign n1293 = ~n1286 & ~n1288;
  assign n1294 = ~n1290 & n1293;
  assign n1295 = ~n1292 & n1294;
  assign 7604 = 137 & ~n1295;
  assign n1297 = ~577 & ~7363;
  assign n1298 = ~580 & n1297;
  assign n1299 = 577 & ~7473;
  assign n1300 = ~580 & n1299;
  assign n1301 = 188 & ~577;
  assign n1302 = 580 & n1301;
  assign n1303 = 158 & 577;
  assign n1304 = 580 & n1303;
  assign n1305 = ~n1298 & ~n1300;
  assign n1306 = ~n1302 & n1305;
  assign n1307 = ~n1304 & n1306;
  assign 7605 = 137 & ~n1307;
  assign n1309 = ~577 & ~7467;
  assign n1310 = ~580 & n1309;
  assign n1311 = 577 & ~7472;
  assign n1312 = ~580 & n1311;
  assign n1313 = 155 & ~577;
  assign n1314 = 580 & n1313;
  assign n1315 = 152 & 577;
  assign n1316 = 580 & n1315;
  assign n1317 = ~n1310 & ~n1312;
  assign n1318 = ~n1314 & n1317;
  assign n1319 = ~n1316 & n1318;
  assign 7606 = 137 & ~n1319;
  assign n1321 = ~577 & ~7466;
  assign n1322 = ~580 & n1321;
  assign n1323 = 577 & ~7471;
  assign n1324 = ~580 & n1323;
  assign n1325 = 149 & ~577;
  assign n1326 = 580 & n1325;
  assign n1327 = 146 & 577;
  assign n1328 = 580 & n1327;
  assign n1329 = ~n1322 & ~n1324;
  assign n1330 = ~n1326 & n1329;
  assign n1331 = ~n1328 & n1330;
  assign 7607 = 137 & ~n1331;
  assign n1333 = 135 & 631;
  assign n1334 = ~603 & ~n381;
  assign n1335 = ~599 & n1334;
  assign n1336 = 132 & n603;
  assign n1337 = n603 & ~n1336;
  assign n1338 = 132 & ~n1336;
  assign n1339 = ~n1337 & ~n1338;
  assign n1340 = 603 & ~n1339;
  assign n1341 = ~599 & n1340;
  assign n1342 = 123 & ~603;
  assign n1343 = 599 & n1342;
  assign n1344 = 603 & ~7432;
  assign n1345 = 599 & n1344;
  assign n1346 = ~n1335 & ~n1341;
  assign n1347 = ~n1343 & n1346;
  assign n1348 = ~n1345 & n1347;
  assign 7626 = ~n1333 & ~n1348;
  assign n1350 = ~7432 & ~n1339;
  assign n1351 = ~n1339 & ~n1350;
  assign n1352 = ~7432 & ~n1350;
  assign 7698 = n1351 | n1352;
  assign n1354 = ~619 & ~n381;
  assign n1355 = ~625 & n1354;
  assign n1356 = 619 & ~7432;
  assign n1357 = ~625 & n1356;
  assign n1358 = 123 & ~619;
  assign n1359 = 625 & n1358;
  assign n1360 = ~n1355 & ~n1357;
  assign 7699 = ~n1359 & n1360;
  assign n1362 = ~619 & n378;
  assign n1363 = ~625 & n1362;
  assign n1364 = 619 & ~n1116;
  assign n1365 = ~625 & n1364;
  assign n1366 = 121 & ~619;
  assign n1367 = 625 & n1366;
  assign n1368 = ~n1363 & ~n1365;
  assign 7700 = ~n1367 & n1368;
  assign n1370 = ~619 & n375;
  assign n1371 = ~625 & n1370;
  assign n1372 = 619 & ~n1105;
  assign n1373 = ~625 & n1372;
  assign n1374 = 116 & ~619;
  assign n1375 = 625 & n1374;
  assign n1376 = ~n1371 & ~n1373;
  assign 7701 = ~n1375 & n1376;
  assign n1378 = ~619 & n365;
  assign n1379 = ~625 & n1378;
  assign n1380 = 619 & ~n1095;
  assign n1381 = ~625 & n1380;
  assign n1382 = 112 & ~619;
  assign n1383 = 625 & n1382;
  assign n1384 = ~n1379 & ~n1381;
  assign 7702 = ~n1383 & n1384;
  assign n1386 = 386 & 559;
  assign n1387 = 556 & n1386;
  assign n1388 = 552 & n1387;
  assign n1389 = 562 & ~7474;
  assign n1390 = ~7476 & n1389;
  assign n1391 = ~6716 & n1390;
  assign n1392 = ~6877 & n1391;
  assign n1393 = n1388 & n1392;
  assign 7703 = 245 & n1393;
  assign n1395 = ~619 & n521;
  assign n1396 = ~625 & n1395;
  assign n1397 = 619 & ~n1084;
  assign n1398 = ~625 & n1397;
  assign n1399 = 115 & ~619;
  assign n1400 = 625 & n1399;
  assign n1401 = ~n1396 & ~n1398;
  assign 7704 = ~n1400 & n1401;
  assign n1403 = ~619 & n465;
  assign n1404 = ~625 & n1403;
  assign n1405 = 619 & ~n1070;
  assign n1406 = ~625 & n1405;
  assign n1407 = 114 & ~619;
  assign n1408 = 625 & n1407;
  assign n1409 = ~n1404 & ~n1406;
  assign 7705 = ~n1408 & n1409;
  assign n1411 = ~619 & n455;
  assign n1412 = ~625 & n1411;
  assign n1413 = 619 & ~n1058;
  assign n1414 = ~625 & n1413;
  assign n1415 = 53 & ~619;
  assign n1416 = 625 & n1415;
  assign n1417 = ~n1412 & ~n1414;
  assign 7706 = ~n1416 & n1417;
  assign n1419 = ~619 & n445;
  assign n1420 = ~625 & n1419;
  assign n1421 = 619 & ~n1048;
  assign n1422 = ~625 & n1421;
  assign n1423 = 113 & ~619;
  assign n1424 = 625 & n1423;
  assign n1425 = ~n1420 & ~n1422;
  assign 7707 = ~n1424 & n1425;
  assign n1427 = ~613 & ~7699;
  assign n1428 = ~616 & n1427;
  assign n1429 = 613 & ~7704;
  assign n1430 = ~616 & n1429;
  assign n1431 = 109 & ~613;
  assign n1432 = 616 & n1431;
  assign n1433 = 106 & 613;
  assign n1434 = 616 & n1433;
  assign n1435 = ~n1428 & ~n1430;
  assign n1436 = ~n1432 & n1435;
  assign 7735 = n1434 | ~n1436;
  assign n1438 = ~610 & ~7699;
  assign n1439 = ~607 & n1438;
  assign n1440 = 610 & ~7704;
  assign n1441 = ~607 & n1440;
  assign n1442 = 109 & ~610;
  assign n1443 = 607 & n1442;
  assign n1444 = 106 & 610;
  assign n1445 = 607 & n1444;
  assign n1446 = ~n1439 & ~n1441;
  assign n1447 = ~n1443 & n1446;
  assign 7736 = n1445 | ~n1447;
  assign n1449 = ~610 & ~7700;
  assign n1450 = ~607 & n1449;
  assign n1451 = 610 & ~7705;
  assign n1452 = ~607 & n1451;
  assign n1453 = 46 & ~610;
  assign n1454 = 607 & n1453;
  assign n1455 = 49 & 610;
  assign n1456 = 607 & n1455;
  assign n1457 = ~n1450 & ~n1452;
  assign n1458 = ~n1454 & n1457;
  assign 7737 = n1456 | ~n1458;
  assign n1460 = ~610 & ~7701;
  assign n1461 = ~607 & n1460;
  assign n1462 = 610 & ~7706;
  assign n1463 = ~607 & n1462;
  assign n1464 = 100 & ~610;
  assign n1465 = 607 & n1464;
  assign n1466 = 103 & 610;
  assign n1467 = 607 & n1466;
  assign n1468 = ~n1461 & ~n1463;
  assign n1469 = ~n1465 & n1468;
  assign 7738 = n1467 | ~n1469;
  assign n1471 = ~610 & ~7702;
  assign n1472 = ~607 & n1471;
  assign n1473 = 610 & ~7707;
  assign n1474 = ~607 & n1473;
  assign n1475 = 91 & ~610;
  assign n1476 = 607 & n1475;
  assign n1477 = 40 & 610;
  assign n1478 = 607 & n1477;
  assign n1479 = ~n1472 & ~n1474;
  assign n1480 = ~n1476 & n1479;
  assign 7739 = n1478 | ~n1480;
  assign n1482 = ~613 & ~7700;
  assign n1483 = ~616 & n1482;
  assign n1484 = 613 & ~7705;
  assign n1485 = ~616 & n1484;
  assign n1486 = 46 & ~613;
  assign n1487 = 616 & n1486;
  assign n1488 = 49 & 613;
  assign n1489 = 616 & n1488;
  assign n1490 = ~n1483 & ~n1485;
  assign n1491 = ~n1487 & n1490;
  assign 7740 = n1489 | ~n1491;
  assign n1493 = ~613 & ~7701;
  assign n1494 = ~616 & n1493;
  assign n1495 = 613 & ~7706;
  assign n1496 = ~616 & n1495;
  assign n1497 = 100 & ~613;
  assign n1498 = 616 & n1497;
  assign n1499 = 103 & 613;
  assign n1500 = 616 & n1499;
  assign n1501 = ~n1494 & ~n1496;
  assign n1502 = ~n1498 & n1501;
  assign 7741 = n1500 | ~n1502;
  assign n1504 = ~613 & ~7702;
  assign n1505 = ~616 & n1504;
  assign n1506 = 613 & ~7707;
  assign n1507 = ~616 & n1506;
  assign n1508 = 91 & ~613;
  assign n1509 = 616 & n1508;
  assign n1510 = 40 & 613;
  assign n1511 = 616 & n1510;
  assign n1512 = ~n1505 & ~n1507;
  assign n1513 = ~n1509 & n1512;
  assign 7742 = n1511 | ~n1513;
  assign n1515 = ~571 & ~7702;
  assign n1516 = ~574 & n1515;
  assign n1517 = 571 & ~7707;
  assign n1518 = ~574 & n1517;
  assign n1519 = 203 & ~571;
  assign n1520 = 574 & n1519;
  assign n1521 = 173 & 571;
  assign n1522 = 574 & n1521;
  assign n1523 = ~n1516 & ~n1518;
  assign n1524 = ~n1520 & n1523;
  assign n1525 = ~n1522 & n1524;
  assign 7754 = 137 & ~n1525;
  assign n1527 = ~571 & ~7701;
  assign n1528 = ~574 & n1527;
  assign n1529 = 571 & ~7706;
  assign n1530 = ~574 & n1529;
  assign n1531 = 197 & ~571;
  assign n1532 = 574 & n1531;
  assign n1533 = 167 & 571;
  assign n1534 = 574 & n1533;
  assign n1535 = ~n1528 & ~n1530;
  assign n1536 = ~n1532 & n1535;
  assign n1537 = ~n1534 & n1536;
  assign 7755 = 137 & ~n1537;
  assign n1539 = ~571 & ~7700;
  assign n1540 = ~574 & n1539;
  assign n1541 = 571 & ~7705;
  assign n1542 = ~574 & n1541;
  assign n1543 = 194 & ~571;
  assign n1544 = 574 & n1543;
  assign n1545 = 164 & 571;
  assign n1546 = 574 & n1545;
  assign n1547 = ~n1540 & ~n1542;
  assign n1548 = ~n1544 & n1547;
  assign n1549 = ~n1546 & n1548;
  assign 7756 = 137 & ~n1549;
  assign n1551 = ~571 & ~7699;
  assign n1552 = ~574 & n1551;
  assign n1553 = 571 & ~7704;
  assign n1554 = ~574 & n1553;
  assign n1555 = 191 & ~571;
  assign n1556 = 574 & n1555;
  assign n1557 = 161 & 571;
  assign n1558 = 574 & n1557;
  assign n1559 = ~n1552 & ~n1554;
  assign n1560 = ~n1556 & n1559;
  assign n1561 = ~n1558 & n1560;
  assign 7757 = 137 & ~n1561;
  assign n1563 = ~577 & ~7702;
  assign n1564 = ~580 & n1563;
  assign n1565 = 577 & ~7707;
  assign n1566 = ~580 & n1565;
  assign n1567 = 203 & ~577;
  assign n1568 = 580 & n1567;
  assign n1569 = 173 & 577;
  assign n1570 = 580 & n1569;
  assign n1571 = ~n1564 & ~n1566;
  assign n1572 = ~n1568 & n1571;
  assign n1573 = ~n1570 & n1572;
  assign 7758 = 137 & ~n1573;
  assign n1575 = ~577 & ~7701;
  assign n1576 = ~580 & n1575;
  assign n1577 = 577 & ~7706;
  assign n1578 = ~580 & n1577;
  assign n1579 = 197 & ~577;
  assign n1580 = 580 & n1579;
  assign n1581 = 167 & 577;
  assign n1582 = 580 & n1581;
  assign n1583 = ~n1576 & ~n1578;
  assign n1584 = ~n1580 & n1583;
  assign n1585 = ~n1582 & n1584;
  assign 7759 = 137 & ~n1585;
  assign n1587 = ~577 & ~7700;
  assign n1588 = ~580 & n1587;
  assign n1589 = 577 & ~7705;
  assign n1590 = ~580 & n1589;
  assign n1591 = 194 & ~577;
  assign n1592 = 580 & n1591;
  assign n1593 = 164 & 577;
  assign n1594 = 580 & n1593;
  assign n1595 = ~n1588 & ~n1590;
  assign n1596 = ~n1592 & n1595;
  assign n1597 = ~n1594 & n1596;
  assign 7760 = 137 & ~n1597;
  assign n1599 = ~577 & ~7699;
  assign n1600 = ~580 & n1599;
  assign n1601 = 577 & ~7704;
  assign n1602 = ~580 & n1601;
  assign n1603 = 191 & ~577;
  assign n1604 = 580 & n1603;
  assign n1605 = 161 & 577;
  assign n1606 = 580 & n1605;
  assign n1607 = ~n1600 & ~n1602;
  assign n1608 = ~n1604 & n1607;
  assign n1609 = ~n1606 & n1608;
  assign 7761 = 137 & ~n1609;
  assign n1611 = n365 & ~n375;
  assign n1612 = ~n365 & n375;
  assign n1613 = ~n1611 & ~n1612;
  assign n1614 = n378 & n381;
  assign n1615 = ~n378 & ~n381;
  assign n1616 = ~n1614 & ~n1615;
  assign n1617 = ~n1613 & n1616;
  assign n1618 = n1613 & ~n1616;
  assign n1619 = ~n1617 & ~n1618;
  assign n1620 = 248 & 534;
  assign n1621 = 351 & n1620;
  assign n1622 = 251 & 534;
  assign n1623 = ~351 & n1622;
  assign n1624 = ~n1621 & ~n1623;
  assign n1625 = 242 & 351;
  assign n1626 = 254 & ~351;
  assign n1627 = ~n1625 & ~n1626;
  assign n1628 = ~534 & n1627;
  assign n1629 = n1624 & ~n1628;
  assign n1630 = 248 & 523;
  assign n1631 = 341 & n1630;
  assign n1632 = 251 & 523;
  assign n1633 = ~341 & n1632;
  assign n1634 = ~n1631 & ~n1633;
  assign n1635 = 242 & 341;
  assign n1636 = 254 & ~341;
  assign n1637 = ~n1635 & ~n1636;
  assign n1638 = ~523 & n1637;
  assign n1639 = n1634 & ~n1638;
  assign n1640 = n1629 & ~n1639;
  assign n1641 = ~n1629 & n1639;
  assign n1642 = ~n1640 & ~n1641;
  assign n1643 = 248 & 514;
  assign n1644 = ~242 & ~514;
  assign n1645 = ~n1643 & ~n1644;
  assign n1646 = 248 & 503;
  assign n1647 = 324 & n1646;
  assign n1648 = 251 & 503;
  assign n1649 = ~324 & n1648;
  assign n1650 = ~n1647 & ~n1649;
  assign n1651 = 242 & 324;
  assign n1652 = 254 & ~324;
  assign n1653 = ~n1651 & ~n1652;
  assign n1654 = ~503 & n1653;
  assign n1655 = n1650 & ~n1654;
  assign n1656 = n1645 & ~n1655;
  assign n1657 = ~n1645 & n1655;
  assign n1658 = ~n1656 & ~n1657;
  assign n1659 = ~n423 & n1642;
  assign n1660 = n1658 & n1659;
  assign n1661 = n423 & n1642;
  assign n1662 = ~n1658 & n1661;
  assign n1663 = ~n1660 & ~n1662;
  assign n1664 = n423 & ~n1642;
  assign n1665 = n1658 & n1664;
  assign n1666 = ~n423 & ~n1642;
  assign n1667 = ~n1658 & n1666;
  assign n1668 = ~n1665 & ~n1667;
  assign n1669 = n1663 & n1668;
  assign n1670 = ~n1619 & n1669;
  assign n1671 = n1619 & ~n1669;
  assign n1672 = ~n1670 & ~n1671;
  assign n1673 = ~619 & n1672;
  assign n1674 = ~625 & n1673;
  assign n1675 = n614 & n873;
  assign n1676 = ~n614 & ~n873;
  assign n1677 = ~n1675 & ~n1676;
  assign n1678 = n888 & n1677;
  assign n1679 = ~n888 & ~n1677;
  assign n1680 = ~n1678 & ~n1679;
  assign n1681 = n859 & n1680;
  assign n1682 = ~n859 & ~n1680;
  assign n1683 = ~n1681 & ~n1682;
  assign n1684 = n614 & n1683;
  assign n1685 = ~n614 & ~n1683;
  assign n1686 = ~n1684 & ~n1685;
  assign n1687 = ~n632 & n1686;
  assign n1688 = n632 & ~n1686;
  assign n1689 = ~n1687 & ~n1688;
  assign n1690 = ~n626 & n1689;
  assign n1691 = n626 & ~n1689;
  assign n1692 = ~n1690 & ~n1691;
  assign n1693 = ~n620 & n1692;
  assign n1694 = n620 & ~n1692;
  assign n1695 = ~n1693 & ~n1694;
  assign n1696 = ~n611 & n1695;
  assign n1697 = n611 & ~n1695;
  assign n1698 = ~n1696 & ~n1697;
  assign n1699 = ~583 & n1698;
  assign n1700 = n614 & ~n620;
  assign n1701 = ~n611 & n1700;
  assign n1702 = ~n632 & n1701;
  assign n1703 = n859 & ~n1702;
  assign n1704 = ~n641 & n888;
  assign n1705 = ~n632 & n1700;
  assign n1706 = n873 & ~n1705;
  assign n1707 = ~n1704 & n1706;
  assign n1708 = n1704 & ~n1706;
  assign n1709 = ~n1707 & ~n1708;
  assign n1710 = ~n1703 & n1709;
  assign n1711 = n1703 & ~n1709;
  assign n1712 = ~n1710 & ~n1711;
  assign n1713 = n614 & n1712;
  assign n1714 = ~n614 & ~n1712;
  assign n1715 = ~n1713 & ~n1714;
  assign n1716 = ~n632 & n1715;
  assign n1717 = n632 & ~n1715;
  assign n1718 = ~n1716 & ~n1717;
  assign n1719 = ~n626 & n1718;
  assign n1720 = n626 & ~n1718;
  assign n1721 = ~n1719 & ~n1720;
  assign n1722 = ~n620 & n1721;
  assign n1723 = n620 & ~n1721;
  assign n1724 = ~n1722 & ~n1723;
  assign n1725 = ~n611 & n1724;
  assign n1726 = n611 & ~n1724;
  assign n1727 = ~n1725 & ~n1726;
  assign n1728 = 583 & ~n1727;
  assign n1729 = ~n1699 & ~n1728;
  assign n1730 = ~n753 & n1106;
  assign n1731 = n753 & ~n1106;
  assign n1732 = ~n1730 & ~n1731;
  assign n1733 = n823 & n1732;
  assign n1734 = ~n823 & ~n1732;
  assign n1735 = ~n1733 & ~n1734;
  assign n1736 = ~n594 & n1735;
  assign n1737 = n594 & ~n1735;
  assign n1738 = ~n1736 & ~n1737;
  assign n1739 = ~n600 & n1738;
  assign n1740 = n600 & ~n1738;
  assign n1741 = ~n1739 & ~n1740;
  assign n1742 = n603 & n1741;
  assign n1743 = ~n603 & ~n1741;
  assign n1744 = ~n1742 & ~n1743;
  assign n1745 = n588 & n1744;
  assign n1746 = ~n588 & ~n1744;
  assign n1747 = ~n1745 & ~n1746;
  assign n1748 = n777 & ~n1747;
  assign n1749 = ~583 & n1748;
  assign n1750 = ~n1100 & ~n1111;
  assign n1751 = n1100 & n1111;
  assign n1752 = ~n1750 & ~n1751;
  assign n1753 = ~n830 & n1752;
  assign n1754 = n830 & ~n1752;
  assign n1755 = ~n1753 & ~n1754;
  assign n1756 = ~n594 & n1755;
  assign n1757 = n594 & ~n1755;
  assign n1758 = ~n1756 & ~n1757;
  assign n1759 = ~n600 & n1758;
  assign n1760 = n600 & ~n1758;
  assign n1761 = ~n1759 & ~n1760;
  assign n1762 = n603 & n1761;
  assign n1763 = ~n603 & ~n1761;
  assign n1764 = ~n1762 & ~n1763;
  assign n1765 = n588 & n1764;
  assign n1766 = ~n588 & ~n1764;
  assign n1767 = ~n1765 & ~n1766;
  assign n1768 = ~n777 & ~n1767;
  assign n1769 = ~583 & n1768;
  assign n1770 = ~n644 & n777;
  assign n1771 = ~n1747 & n1770;
  assign n1772 = 583 & n1771;
  assign n1773 = ~n1767 & ~n1770;
  assign n1774 = 583 & n1773;
  assign n1775 = ~n1749 & ~n1769;
  assign n1776 = ~n1772 & n1775;
  assign n1777 = ~n1774 & n1776;
  assign n1778 = ~n1729 & n1777;
  assign n1779 = n1729 & ~n1777;
  assign n1780 = ~n1778 & ~n1779;
  assign n1781 = 619 & ~n1780;
  assign n1782 = ~625 & n1781;
  assign n1783 = 120 & ~619;
  assign n1784 = 625 & n1783;
  assign n1785 = 619 & 625;
  assign n1786 = ~n1674 & ~n1782;
  assign n1787 = ~n1784 & n1786;
  assign 8075 = n1785 | ~n1787;
  assign n1789 = 248 & 422;
  assign n1790 = 226 & n1789;
  assign n1791 = 251 & 422;
  assign n1792 = ~226 & n1791;
  assign n1793 = ~n1790 & ~n1792;
  assign n1794 = 226 & 242;
  assign n1795 = ~226 & 254;
  assign n1796 = ~n1794 & ~n1795;
  assign n1797 = ~422 & n1796;
  assign n1798 = n1793 & ~n1797;
  assign n1799 = 248 & 468;
  assign n1800 = 218 & n1799;
  assign n1801 = 251 & 468;
  assign n1802 = ~218 & n1801;
  assign n1803 = ~n1800 & ~n1802;
  assign n1804 = 218 & 242;
  assign n1805 = ~218 & 254;
  assign n1806 = ~n1804 & ~n1805;
  assign n1807 = ~468 & n1806;
  assign n1808 = n1803 & ~n1807;
  assign n1809 = n1798 & ~n1808;
  assign n1810 = ~n1798 & n1808;
  assign n1811 = ~n1809 & ~n1810;
  assign n1812 = 248 & 457;
  assign n1813 = 210 & n1812;
  assign n1814 = 251 & 457;
  assign n1815 = ~210 & n1814;
  assign n1816 = ~n1813 & ~n1815;
  assign n1817 = 210 & 242;
  assign n1818 = ~210 & 254;
  assign n1819 = ~n1817 & ~n1818;
  assign n1820 = ~457 & n1819;
  assign n1821 = n1816 & ~n1820;
  assign n1822 = ~n521 & n1821;
  assign n1823 = n521 & ~n1821;
  assign n1824 = ~n1822 & ~n1823;
  assign n1825 = ~n1811 & n1824;
  assign n1826 = n1811 & ~n1824;
  assign n1827 = ~n1825 & ~n1826;
  assign n1828 = 248 & 374;
  assign n1829 = 281 & n1828;
  assign n1830 = 251 & 374;
  assign n1831 = ~281 & n1830;
  assign n1832 = ~n1829 & ~n1831;
  assign n1833 = 242 & 281;
  assign n1834 = 254 & ~281;
  assign n1835 = ~n1833 & ~n1834;
  assign n1836 = ~374 & n1835;
  assign n1837 = n1832 & ~n1836;
  assign n1838 = 248 & 411;
  assign n1839 = 273 & n1838;
  assign n1840 = 251 & 411;
  assign n1841 = ~273 & n1840;
  assign n1842 = ~n1839 & ~n1841;
  assign n1843 = 242 & 273;
  assign n1844 = 254 & ~273;
  assign n1845 = ~n1843 & ~n1844;
  assign n1846 = ~411 & n1845;
  assign n1847 = n1842 & ~n1846;
  assign n1848 = 248 & 400;
  assign n1849 = 265 & n1848;
  assign n1850 = 251 & 400;
  assign n1851 = ~265 & n1850;
  assign n1852 = ~n1849 & ~n1851;
  assign n1853 = 242 & 265;
  assign n1854 = 254 & ~265;
  assign n1855 = ~n1853 & ~n1854;
  assign n1856 = ~400 & n1855;
  assign n1857 = n1852 & ~n1856;
  assign n1858 = n1847 & ~n1857;
  assign n1859 = ~n1847 & n1857;
  assign n1860 = ~n1858 & ~n1859;
  assign n1861 = 248 & 389;
  assign n1862 = 257 & n1861;
  assign n1863 = 251 & 389;
  assign n1864 = ~257 & n1863;
  assign n1865 = ~n1862 & ~n1864;
  assign n1866 = 242 & 257;
  assign n1867 = 254 & ~257;
  assign n1868 = ~n1866 & ~n1867;
  assign n1869 = ~389 & n1868;
  assign n1870 = n1865 & ~n1869;
  assign n1871 = 248 & 435;
  assign n1872 = 234 & n1871;
  assign n1873 = 251 & 435;
  assign n1874 = ~234 & n1873;
  assign n1875 = ~n1872 & ~n1874;
  assign n1876 = 234 & 242;
  assign n1877 = ~234 & 254;
  assign n1878 = ~n1876 & ~n1877;
  assign n1879 = ~435 & n1878;
  assign n1880 = n1875 & ~n1879;
  assign n1881 = n1870 & ~n1880;
  assign n1882 = ~n1870 & n1880;
  assign n1883 = ~n1881 & ~n1882;
  assign n1884 = ~n1837 & n1860;
  assign n1885 = n1883 & n1884;
  assign n1886 = n1837 & n1860;
  assign n1887 = ~n1883 & n1886;
  assign n1888 = ~n1885 & ~n1887;
  assign n1889 = n1837 & ~n1860;
  assign n1890 = n1883 & n1889;
  assign n1891 = ~n1837 & ~n1860;
  assign n1892 = ~n1883 & n1891;
  assign n1893 = ~n1890 & ~n1892;
  assign n1894 = n1888 & n1893;
  assign n1895 = ~n1827 & n1894;
  assign n1896 = n1827 & ~n1894;
  assign n1897 = ~n1895 & ~n1896;
  assign n1898 = ~619 & n1897;
  assign n1899 = ~625 & n1898;
  assign n1900 = ~n738 & n937;
  assign n1901 = n738 & ~n937;
  assign n1902 = ~n1900 & ~n1901;
  assign n1903 = n952 & n1902;
  assign n1904 = ~n952 & ~n1902;
  assign n1905 = ~n1903 & ~n1904;
  assign n1906 = n923 & n1905;
  assign n1907 = ~n923 & ~n1905;
  assign n1908 = ~n1906 & ~n1907;
  assign n1909 = ~n556 & n1908;
  assign n1910 = n556 & ~n1908;
  assign n1911 = ~n1909 & ~n1910;
  assign n1912 = ~n562 & n1911;
  assign n1913 = n562 & ~n1911;
  assign n1914 = ~n1912 & ~n1913;
  assign n1915 = ~n580 & n1914;
  assign n1916 = n580 & ~n1914;
  assign n1917 = ~n1915 & ~n1916;
  assign n1918 = ~n568 & n1917;
  assign n1919 = n568 & ~n1917;
  assign n1920 = ~n1918 & ~n1919;
  assign n1921 = ~n574 & n1920;
  assign n1922 = n574 & ~n1920;
  assign n1923 = ~n1921 & ~n1922;
  assign n1924 = ~566 & n1923;
  assign n1925 = ~n556 & ~n568;
  assign n1926 = ~n574 & n1925;
  assign n1927 = ~n562 & n1926;
  assign n1928 = n923 & ~n1927;
  assign n1929 = ~n581 & n952;
  assign n1930 = ~n562 & n1925;
  assign n1931 = n937 & ~n1930;
  assign n1932 = ~374 & n553;
  assign n1933 = ~n1931 & ~n1932;
  assign n1934 = n1931 & n1932;
  assign n1935 = ~n1933 & ~n1934;
  assign n1936 = ~n1929 & n1935;
  assign n1937 = n1929 & ~n1935;
  assign n1938 = ~n1936 & ~n1937;
  assign n1939 = ~n1928 & n1938;
  assign n1940 = n1928 & ~n1938;
  assign n1941 = ~n1939 & ~n1940;
  assign n1942 = ~n556 & n1941;
  assign n1943 = n556 & ~n1941;
  assign n1944 = ~n1942 & ~n1943;
  assign n1945 = ~n562 & n1944;
  assign n1946 = n562 & ~n1944;
  assign n1947 = ~n1945 & ~n1946;
  assign n1948 = ~n580 & n1947;
  assign n1949 = n580 & ~n1947;
  assign n1950 = ~n1948 & ~n1949;
  assign n1951 = ~n568 & n1950;
  assign n1952 = n568 & ~n1950;
  assign n1953 = ~n1951 & ~n1952;
  assign n1954 = ~n574 & n1953;
  assign n1955 = n574 & ~n1953;
  assign n1956 = ~n1954 & ~n1955;
  assign n1957 = 566 & ~n1956;
  assign n1958 = ~n1924 & ~n1957;
  assign n1959 = ~n721 & n1060;
  assign n1960 = n721 & ~n1060;
  assign n1961 = ~n1959 & ~n1960;
  assign n1962 = n1074 & n1961;
  assign n1963 = ~n1074 & ~n1961;
  assign n1964 = ~n1962 & ~n1963;
  assign n1965 = ~n529 & n1964;
  assign n1966 = n529 & ~n1964;
  assign n1967 = ~n1965 & ~n1966;
  assign n1968 = ~n535 & n1967;
  assign n1969 = n535 & ~n1967;
  assign n1970 = ~n1968 & ~n1969;
  assign n1971 = ~n547 & n1970;
  assign n1972 = n547 & ~n1970;
  assign n1973 = ~n1971 & ~n1972;
  assign n1974 = ~n541 & n1973;
  assign n1975 = n541 & ~n1973;
  assign n1976 = ~n1974 & ~n1975;
  assign n1977 = n746 & ~n1976;
  assign n1978 = ~566 & n1977;
  assign n1979 = ~n1053 & ~n1065;
  assign n1980 = n1053 & n1065;
  assign n1981 = ~n1979 & ~n1980;
  assign n1982 = ~n1079 & n1981;
  assign n1983 = n1079 & ~n1981;
  assign n1984 = ~n1982 & ~n1983;
  assign n1985 = ~n529 & n1984;
  assign n1986 = n529 & ~n1984;
  assign n1987 = ~n1985 & ~n1986;
  assign n1988 = ~n535 & n1987;
  assign n1989 = n535 & ~n1987;
  assign n1990 = ~n1988 & ~n1989;
  assign n1991 = ~n547 & n1990;
  assign n1992 = n547 & ~n1990;
  assign n1993 = ~n1991 & ~n1992;
  assign n1994 = ~n541 & n1993;
  assign n1995 = n541 & ~n1993;
  assign n1996 = ~n1994 & ~n1995;
  assign n1997 = ~n746 & ~n1996;
  assign n1998 = ~566 & n1997;
  assign n1999 = ~n584 & n746;
  assign n2000 = ~n1976 & n1999;
  assign n2001 = 566 & n2000;
  assign n2002 = ~n1996 & ~n1999;
  assign n2003 = 566 & n2002;
  assign n2004 = ~n1978 & ~n1998;
  assign n2005 = ~n2001 & n2004;
  assign n2006 = ~n2003 & n2005;
  assign n2007 = ~n1958 & n2006;
  assign n2008 = n1958 & ~n2006;
  assign n2009 = ~n2007 & ~n2008;
  assign n2010 = 619 & ~n2009;
  assign n2011 = ~625 & n2010;
  assign n2012 = 118 & ~619;
  assign n2013 = 625 & n2012;
  assign n2014 = ~n1899 & ~n2011;
  assign n2015 = ~n2013 & n2014;
  assign 8076 = n1785 | ~n2015;
  assign n2017 = ~619 & ~n1672;
  assign n2018 = 619 & n1780;
  assign n2019 = ~n2017 & ~n2018;
  assign n2020 = ~625 & ~n2019;
  assign n2021 = 94 & 625;
  assign n2022 = ~n2020 & ~n2021;
  assign n2023 = ~610 & ~n2022;
  assign n2024 = ~607 & n2023;
  assign n2025 = ~619 & ~n1897;
  assign n2026 = 619 & n2009;
  assign n2027 = ~n2025 & ~n2026;
  assign n2028 = ~625 & ~n2027;
  assign n2029 = 97 & 625;
  assign n2030 = ~n2028 & ~n2029;
  assign n2031 = 610 & ~n2030;
  assign n2032 = ~607 & n2031;
  assign n2033 = 14 & ~610;
  assign n2034 = 607 & n2033;
  assign n2035 = 64 & 610;
  assign n2036 = 607 & n2035;
  assign n2037 = ~n2024 & ~n2032;
  assign n2038 = ~n2034 & n2037;
  assign 8123 = n2036 | ~n2038;
  assign n2040 = ~613 & ~n2022;
  assign n2041 = ~616 & n2040;
  assign n2042 = 613 & ~n2030;
  assign n2043 = ~616 & n2042;
  assign n2044 = 14 & ~613;
  assign n2045 = 616 & n2044;
  assign n2046 = 64 & 613;
  assign n2047 = 616 & n2046;
  assign n2048 = ~n2041 & ~n2043;
  assign n2049 = ~n2045 & n2048;
  assign 8124 = n2047 | ~n2049;
  assign n2051 = ~571 & ~n2022;
  assign n2052 = ~574 & n2051;
  assign n2053 = 571 & ~n2030;
  assign n2054 = ~574 & n2053;
  assign n2055 = 176 & ~571;
  assign n2056 = 574 & n2055;
  assign n2057 = 179 & 571;
  assign n2058 = 574 & n2057;
  assign n2059 = ~n2052 & ~n2054;
  assign n2060 = ~n2056 & n2059;
  assign n2061 = ~n2058 & n2060;
  assign 8127 = ~137 | n2061;
  assign n2063 = ~577 & ~n2022;
  assign n2064 = ~580 & n2063;
  assign n2065 = 577 & ~n2030;
  assign n2066 = ~580 & n2065;
  assign n2067 = 176 & ~577;
  assign n2068 = 580 & n2067;
  assign n2069 = 179 & 577;
  assign n2070 = 580 & n2069;
  assign n2071 = ~n2064 & ~n2066;
  assign n2072 = ~n2068 & n2071;
  assign n2073 = ~n2070 & n2072;
  assign 8128 = ~137 | n2073;
  assign 1137 = ~545;
  assign 1138 = ~348;
  assign 1139 = ~366;
  assign 1141 = ~549;
  assign 1144 = ~338;
  assign 1145 = ~358;
  assign 1152 = ~245;
  assign 1153 = ~552;
  assign 1154 = ~562;
  assign 1155 = ~559;
  assign 3613 = ~299;
  assign 709 = 141;
  assign 816 = 293;
  assign 1066 = 592;
  assign 1142 = 1137;
  assign 1143 = 1137;
  assign 2139 = 137;
  assign 2142 = 141;
  assign 2309 = \1 ;
  assign 2387 = 549;
  assign 2527 = 299;
  assign 2584 = 1141;
  assign 3357 = \1 ;
  assign 3358 = \1 ;
  assign 3359 = \1 ;
  assign 3360 = \1 ;
  assign 3604 = 299;
  assign 4278 = 4275;
endmodule
