module top (
    \1 , 2, 3, 4, 5, 6, 7, 8, 11, 14, 15, 16, 19, 20, 21, 22, 23, 24, 25,
    26, 27, 28, 29, 32, 33, 34, 35, 36, 37, 40, 43, 44, 47, 48, 49, 50, 51,
    52, 53, 54, 55, 56, 57, 60, 61, 62, 63, 64, 65, 66, 67, 68, 69, 72, 73,
    74, 75, 76, 77, 78, 79, 80, 81, 82, 85, 86, 87, 88, 89, 90, 91, 92, 93,
    94, 95, 96, 99, 100, 101, 102, 103, 104, 105, 106, 107, 108, 111, 112,
    113, 114, 115, 116, 117, 118, 119, 120, 123, 124, 125, 126, 127, 128,
    129, 130, 131, 132, 135, 136, 137, 138, 139, 140, 141, 142, 143, 144,
    145, 146, 147, 148, 149, 150, 151, 152, 153, 154, 155, 156, 157, 158,
    159, 160, 161, 162, 163, 164, 165, 166, 167, 168, 169, 170, 171, 172,
    173, 174, 175, 176, 177, 178, 179, 180, 181, 182, 183, 184, 185, 186,
    187, 188, 189, 190, 191, 192, 193, 194, 195, 196, 197, 198, 199, 200,
    201, 202, 203, 204, 205, 206, 207, 208, 209, 210, 211, 212, 213, 214,
    215, 216, 217, 218, 219, 224, 227, 230, 231, 234, 237, 241, 246, 253,
    256, 259, 262, 263, 266, 269, 272, 275, 278, 281, 284, 287, 290, 294,
    297, 301, 305, 309, 313, 316, 319, 322, 325, 328, 331, 334, 337, 340,
    343, 346, 349, 352, 355,
    398, 400, 401, 419, 420, 456, 457, 458, 487, 488, 489, 490, 491, 492,
    493, 494, 792, 799, 805, 1026, 1028, 1029, 1269, 1277, 1448, 1726,
    1816, 1817, 1818, 1819, 1820, 1821, 1969, 1970, 1971, 2010, 2012, 2014,
    2016, 2018, 2020, 2022, 2387, 2388, 2389, 2390, 2496, 2643, 2644, 2891,
    2925, 2970, 2971, 3038, 3079, 3546, 3671, 3803, 3804, 3809, 3851, 3875,
    3881, 3882  );
  input  \1 , 2, 3, 4, 5, 6, 7, 8, 11, 14, 15, 16, 19, 20, 21, 22, 23,
    24, 25, 26, 27, 28, 29, 32, 33, 34, 35, 36, 37, 40, 43, 44, 47, 48, 49,
    50, 51, 52, 53, 54, 55, 56, 57, 60, 61, 62, 63, 64, 65, 66, 67, 68, 69,
    72, 73, 74, 75, 76, 77, 78, 79, 80, 81, 82, 85, 86, 87, 88, 89, 90, 91,
    92, 93, 94, 95, 96, 99, 100, 101, 102, 103, 104, 105, 106, 107, 108,
    111, 112, 113, 114, 115, 116, 117, 118, 119, 120, 123, 124, 125, 126,
    127, 128, 129, 130, 131, 132, 135, 136, 137, 138, 139, 140, 141, 142,
    143, 144, 145, 146, 147, 148, 149, 150, 151, 152, 153, 154, 155, 156,
    157, 158, 159, 160, 161, 162, 163, 164, 165, 166, 167, 168, 169, 170,
    171, 172, 173, 174, 175, 176, 177, 178, 179, 180, 181, 182, 183, 184,
    185, 186, 187, 188, 189, 190, 191, 192, 193, 194, 195, 196, 197, 198,
    199, 200, 201, 202, 203, 204, 205, 206, 207, 208, 209, 210, 211, 212,
    213, 214, 215, 216, 217, 218, 219, 224, 227, 230, 231, 234, 237, 241,
    246, 253, 256, 259, 262, 263, 266, 269, 272, 275, 278, 281, 284, 287,
    290, 294, 297, 301, 305, 309, 313, 316, 319, 322, 325, 328, 331, 334,
    337, 340, 343, 346, 349, 352, 355;
  output 398, 400, 401, 419, 420, 456, 457, 458, 487, 488, 489, 490, 491, 492,
    493, 494, 792, 799, 805, 1026, 1028, 1029, 1269, 1277, 1448, 1726,
    1816, 1817, 1818, 1819, 1820, 1821, 1969, 1970, 1971, 2010, 2012, 2014,
    2016, 2018, 2020, 2022, 2387, 2388, 2389, 2390, 2496, 2643, 2644, 2891,
    2925, 2970, 2971, 3038, 3079, 3546, 3671, 3803, 3804, 3809, 3851, 3875,
    3881, 3882;
  wire n375, n376, n378, n384, n385, n386, n387, n388, n389, n391, n392,
    n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n405, n406,
    n407, n408, n409, n410, n411, n412, n413, n414, n416, n417, n418, n419,
    n420, n421, n422, n423, n424, n425, n427, n428, n429, n430, n431, n432,
    n433, n434, n435, n436, n438, n439, n440, n441, n442, n443, n444, n445,
    n446, n447, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
    n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
    n473, n474, n476, n477, n479, n480, n481, n482, n483, n484, n485, n486,
    n487, n488, n490, n491, n492, n493, n494, n495, n496, n497, n498, n500,
    n501, n502, n503, n504, n505, n506, n507, n508, n509, n511, n512, n513,
    n514, n515, n516, n517, n518, n519, n520, n522, n523, n524, n525, n526,
    n527, n528, n529, n530, n531, n532, n533, n534, n536, n537, n539, n540,
    n541, n543, n544, n546, n547, n548, n549, n550, n551, n552, n553, n554,
    n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
    n567, n568, n569, n570, n571, n573, n574, n575, n576, n577, n578, n579,
    n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
    n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
    n604, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
    n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
    n629, n630, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
    n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
    n654, n655, n656, n657, n658, n659, n660, n661, n662, n664, n665, n666,
    n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
    n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
    n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
    n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
    n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
    n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
    n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
    n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
    n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
    n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786,
    n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798,
    n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810,
    n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
    n823, n824, n825, n827, n828, n829, n830, n831, n832, n833, n834, n835,
    n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847,
    n848, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
    n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
    n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
    n885, n886, n887, n888, n889, n890, n891, n892, n894, n895, n896, n897,
    n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909,
    n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921,
    n922, n923, n924, n926, n927, n928, n929, n930, n931, n932, n933, n934,
    n935, n936, n937, n938, n939, n940, n941, n942, n944, n945, n946, n947,
    n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
    n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
    n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
    n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995,
    n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005,
    n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
    n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
    n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035,
    n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045,
    n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055,
    n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065,
    n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075,
    n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085,
    n1087, n1088, n1089, n1090;
  assign n375 = 305 & 309;
  assign n376 = 301 & n375;
  assign 792 = ~297 | ~n376;
  assign n378 = 2 & 15;
  assign 799 = ~237 | ~n378;
  assign 1026 = 94 & 219;
  assign 1028 = ~7 | ~237;
  assign 1029 = ~231 | 1028;
  assign 1269 = ~325 | 1028;
  assign n384 = 57 & 120;
  assign n385 = 108 & n384;
  assign n386 = 69 & n385;
  assign n387 = 82 & 132;
  assign n388 = 96 & n387;
  assign n389 = 44 & n388;
  assign 1277 = n386 & n389;
  assign n391 = 325 & ~n389;
  assign n392 = 231 & ~n386;
  assign 1726 = ~n391 & ~n392;
  assign n394 = 137 & ~319;
  assign n395 = ~322 & n394;
  assign n396 = 101 & 319;
  assign n397 = ~322 & n396;
  assign n398 = 125 & ~319;
  assign n399 = 322 & n398;
  assign n400 = 113 & 319;
  assign n401 = 322 & n400;
  assign n402 = ~n395 & ~n397;
  assign n403 = ~n399 & n402;
  assign 1816 = ~n401 & n403;
  assign n405 = 136 & ~319;
  assign n406 = ~322 & n405;
  assign n407 = 100 & 319;
  assign n408 = ~322 & n407;
  assign n409 = 124 & ~319;
  assign n410 = 322 & n409;
  assign n411 = 112 & 319;
  assign n412 = 322 & n411;
  assign n413 = ~n406 & ~n408;
  assign n414 = ~n410 & n413;
  assign 1817 = ~n412 & n414;
  assign n416 = 138 & ~319;
  assign n417 = ~322 & n416;
  assign n418 = 102 & 319;
  assign n419 = ~322 & n418;
  assign n420 = 126 & ~319;
  assign n421 = 322 & n420;
  assign n422 = 114 & 319;
  assign n423 = 322 & n422;
  assign n424 = ~n417 & ~n419;
  assign n425 = ~n421 & n424;
  assign 1818 = ~n423 & n425;
  assign n427 = 88 & ~227;
  assign n428 = ~234 & n427;
  assign n429 = 50 & 227;
  assign n430 = ~234 & n429;
  assign n431 = 62 & ~227;
  assign n432 = 234 & n431;
  assign n433 = 75 & 227;
  assign n434 = 234 & n433;
  assign n435 = ~n428 & ~n430;
  assign n436 = ~n432 & n435;
  assign 1819 = ~n434 & n436;
  assign n438 = 89 & ~227;
  assign n439 = ~234 & n438;
  assign n440 = 51 & 227;
  assign n441 = ~234 & n440;
  assign n442 = 63 & ~227;
  assign n443 = 234 & n442;
  assign n444 = 76 & 227;
  assign n445 = 234 & n444;
  assign n446 = ~n439 & ~n441;
  assign n447 = ~n443 & n446;
  assign 1820 = ~n445 & n447;
  assign n449 = 90 & ~227;
  assign n450 = ~234 & n449;
  assign n451 = 52 & 227;
  assign n452 = ~234 & n451;
  assign n453 = 64 & ~227;
  assign n454 = 234 & n453;
  assign n455 = 77 & 227;
  assign n456 = 234 & n455;
  assign n457 = ~n450 & ~n452;
  assign n458 = ~n454 & n457;
  assign 1821 = ~n456 & n458;
  assign n460 = 81 & ~227;
  assign n461 = ~234 & n460;
  assign n462 = 43 & 227;
  assign n463 = ~234 & n462;
  assign n464 = 56 & ~227;
  assign n465 = 234 & n464;
  assign n466 = 68 & 227;
  assign n467 = 234 & n466;
  assign n468 = ~n461 & ~n463;
  assign n469 = ~n465 & n468;
  assign n470 = ~n467 & n469;
  assign n471 = 241 & ~n470;
  assign 1969 = ~241 | n471;
  assign n473 = 224 & 237;
  assign n474 = 36 & n473;
  assign 1970 = ~1726 | ~n474;
  assign n476 = \1  & 3;
  assign n477 = 1726 & n473;
  assign 1971 = n476 | ~n477;
  assign n479 = 91 & ~227;
  assign n480 = ~234 & n479;
  assign n481 = 53 & 227;
  assign n482 = ~234 & n481;
  assign n483 = 65 & ~227;
  assign n484 = 234 & n483;
  assign n485 = 78 & 227;
  assign n486 = 234 & n485;
  assign n487 = ~n480 & ~n482;
  assign n488 = ~n484 & n487;
  assign 2010 = n486 | ~n488;
  assign n490 = 87 & ~227;
  assign n491 = ~234 & n490;
  assign n492 = 49 & 227;
  assign n493 = ~234 & n492;
  assign n494 = ~227 & 234;
  assign n495 = 74 & 227;
  assign n496 = 234 & n495;
  assign n497 = ~n491 & ~n493;
  assign n498 = ~n494 & n497;
  assign 2018 = n496 | ~n498;
  assign n500 = 86 & ~227;
  assign n501 = ~234 & n500;
  assign n502 = 48 & 227;
  assign n503 = ~234 & n502;
  assign n504 = 61 & ~227;
  assign n505 = 234 & n504;
  assign n506 = 73 & 227;
  assign n507 = 234 & n506;
  assign n508 = ~n501 & ~n503;
  assign n509 = ~n505 & n508;
  assign 2020 = n507 | ~n509;
  assign n511 = 85 & ~227;
  assign n512 = ~234 & n511;
  assign n513 = 47 & 227;
  assign n514 = ~234 & n513;
  assign n515 = 60 & ~227;
  assign n516 = 234 & n515;
  assign n517 = 72 & 227;
  assign n518 = 234 & n517;
  assign n519 = ~n512 & ~n514;
  assign n520 = ~n516 & n519;
  assign 2022 = n518 | ~n520;
  assign n522 = 92 & ~227;
  assign n523 = ~234 & n522;
  assign n524 = 54 & 227;
  assign n525 = ~234 & n524;
  assign n526 = 66 & ~227;
  assign n527 = 234 & n526;
  assign n528 = 79 & 227;
  assign n529 = 234 & n528;
  assign n530 = ~n523 & ~n525;
  assign n531 = ~n527 & n530;
  assign n532 = ~n529 & n531;
  assign n533 = ~246 & ~n532;
  assign n534 = 246 & ~1821;
  assign 2387 = n533 | n534;
  assign n536 = ~246 & 2010;
  assign n537 = 246 & ~1820;
  assign 2389 = n536 | n537;
  assign n539 = ~230 & n532;
  assign n540 = ~241 & ~n539;
  assign n541 = 241 & ~n532;
  assign 2496 = n540 | n541;
  assign n543 = ~246 & ~n470;
  assign n544 = 246 & ~n539;
  assign 2643 = n543 | n544;
  assign n546 = ~319 & ~322;
  assign n547 = 319 & ~322;
  assign n548 = ~319 & 322;
  assign n549 = 319 & 322;
  assign n550 = ~n546 & ~n547;
  assign n551 = ~n548 & n550;
  assign n552 = ~n549 & n551;
  assign n553 = ~316 & ~n552;
  assign n554 = ~316 & ~n553;
  assign n555 = ~n552 & ~n553;
  assign n556 = ~n554 & ~n555;
  assign n557 = 135 & ~319;
  assign n558 = ~322 & n557;
  assign n559 = 99 & 319;
  assign n560 = ~322 & n559;
  assign n561 = 123 & ~319;
  assign n562 = 322 & n561;
  assign n563 = 111 & 319;
  assign n564 = 322 & n563;
  assign n565 = ~n558 & ~n560;
  assign n566 = ~n562 & n565;
  assign n567 = ~n564 & n566;
  assign n568 = ~313 & ~n567;
  assign n569 = ~313 & ~n568;
  assign n570 = ~n567 & ~n568;
  assign n571 = ~n569 & ~n570;
  assign 2891 = ~n556 | ~n571;
  assign n573 = ~346 & 349;
  assign n574 = 346 & ~349;
  assign n575 = ~n573 & ~n574;
  assign n576 = 256 & ~259;
  assign n577 = ~256 & 259;
  assign n578 = ~n576 & ~n577;
  assign n579 = ~n575 & n578;
  assign n580 = n575 & ~n578;
  assign n581 = ~n579 & ~n580;
  assign n582 = ~328 & 331;
  assign n583 = 328 & ~331;
  assign n584 = ~n582 & ~n583;
  assign n585 = ~334 & 337;
  assign n586 = 334 & ~337;
  assign n587 = ~n585 & ~n586;
  assign n588 = ~340 & 343;
  assign n589 = 340 & ~343;
  assign n590 = ~n588 & ~n589;
  assign n591 = ~n584 & n587;
  assign n592 = n590 & n591;
  assign n593 = n584 & n587;
  assign n594 = ~n590 & n593;
  assign n595 = ~n592 & ~n594;
  assign n596 = n584 & ~n587;
  assign n597 = n590 & n596;
  assign n598 = ~n584 & ~n587;
  assign n599 = ~n590 & n598;
  assign n600 = ~n597 & ~n599;
  assign n601 = n595 & n600;
  assign n602 = ~n581 & n601;
  assign n603 = n581 & ~n601;
  assign n604 = ~n602 & ~n603;
  assign 2925 = 14 & n604;
  assign n606 = 313 & ~316;
  assign n607 = ~313 & 316;
  assign n608 = ~n606 & ~n607;
  assign n609 = ~294 & 355;
  assign n610 = 294 & ~355;
  assign n611 = ~n609 & ~n610;
  assign n612 = 297 & ~301;
  assign n613 = ~297 & 301;
  assign n614 = ~n612 & ~n613;
  assign n615 = 305 & ~309;
  assign n616 = ~305 & 309;
  assign n617 = ~n615 & ~n616;
  assign n618 = ~n611 & n614;
  assign n619 = n617 & n618;
  assign n620 = n611 & n614;
  assign n621 = ~n617 & n620;
  assign n622 = ~n619 & ~n621;
  assign n623 = n611 & ~n614;
  assign n624 = n617 & n623;
  assign n625 = ~n611 & ~n614;
  assign n626 = ~n617 & n625;
  assign n627 = ~n624 & ~n626;
  assign n628 = n622 & n627;
  assign n629 = ~n608 & n628;
  assign n630 = n608 & ~n628;
  assign 2970 = ~n629 & ~n630;
  assign n632 = 278 & ~281;
  assign n633 = ~278 & 281;
  assign n634 = ~n632 & ~n633;
  assign n635 = 284 & ~287;
  assign n636 = ~284 & 287;
  assign n637 = ~n635 & ~n636;
  assign n638 = ~n634 & n637;
  assign n639 = n634 & ~n637;
  assign n640 = ~n638 & ~n639;
  assign n641 = ~263 & 352;
  assign n642 = 263 & ~352;
  assign n643 = ~n641 & ~n642;
  assign n644 = 266 & ~269;
  assign n645 = ~266 & 269;
  assign n646 = ~n644 & ~n645;
  assign n647 = 272 & ~275;
  assign n648 = ~272 & 275;
  assign n649 = ~n647 & ~n648;
  assign n650 = ~n643 & n646;
  assign n651 = n649 & n650;
  assign n652 = n643 & n646;
  assign n653 = ~n649 & n652;
  assign n654 = ~n651 & ~n653;
  assign n655 = n643 & ~n646;
  assign n656 = n649 & n655;
  assign n657 = ~n643 & ~n646;
  assign n658 = ~n649 & n657;
  assign n659 = ~n656 & ~n658;
  assign n660 = n654 & n659;
  assign n661 = ~n640 & n660;
  assign n662 = n640 & ~n660;
  assign 2971 = ~n661 & ~n662;
  assign n664 = 25 & ~29;
  assign n665 = 131 & ~319;
  assign n666 = ~322 & n665;
  assign n667 = 95 & 319;
  assign n668 = ~322 & n667;
  assign n669 = 119 & ~319;
  assign n670 = 322 & n669;
  assign n671 = 107 & 319;
  assign n672 = 322 & n671;
  assign n673 = ~n666 & ~n668;
  assign n674 = ~n670 & n673;
  assign n675 = ~n672 & n674;
  assign n676 = 29 & ~n675;
  assign n677 = ~n664 & ~n676;
  assign n678 = 284 & ~n677;
  assign n679 = ~284 & n677;
  assign n680 = ~n678 & ~n679;
  assign n681 = ~16 & 24;
  assign n682 = 16 & 2022;
  assign n683 = ~n681 & ~n682;
  assign n684 = 281 & ~n683;
  assign n685 = ~281 & n683;
  assign n686 = ~n684 & ~n685;
  assign n687 = 6 & ~16;
  assign n688 = 16 & 2020;
  assign n689 = ~n687 & ~n688;
  assign n690 = 278 & ~n689;
  assign n691 = ~278 & n689;
  assign n692 = ~n690 & ~n691;
  assign n693 = ~16 & 23;
  assign n694 = 16 & 2018;
  assign n695 = ~n693 & ~n694;
  assign n696 = 275 & ~n695;
  assign n697 = ~275 & n695;
  assign n698 = ~n696 & ~n697;
  assign n699 = ~16 & 22;
  assign n700 = 16 & ~1819;
  assign n701 = ~n699 & ~n700;
  assign n702 = 272 & ~n701;
  assign n703 = ~272 & n701;
  assign n704 = ~n702 & ~n703;
  assign n705 = n680 & n686;
  assign n706 = n692 & n705;
  assign n707 = n698 & n706;
  assign n708 = n704 & n707;
  assign n709 = ~16 & 21;
  assign n710 = 16 & ~1820;
  assign n711 = ~n709 & ~n710;
  assign n712 = 269 & ~n711;
  assign n713 = ~269 & n711;
  assign n714 = ~n712 & ~n713;
  assign n715 = 5 & ~16;
  assign n716 = 16 & ~1821;
  assign n717 = ~n715 & ~n716;
  assign n718 = 266 & ~n717;
  assign n719 = ~266 & n717;
  assign n720 = ~n718 & ~n719;
  assign n721 = ~16 & 20;
  assign n722 = 16 & 2010;
  assign n723 = ~n721 & ~n722;
  assign n724 = 263 & ~n723;
  assign n725 = ~263 & n723;
  assign n726 = ~n724 & ~n725;
  assign n727 = 4 & ~16;
  assign n728 = 16 & ~n532;
  assign n729 = ~n727 & ~n728;
  assign n730 = 259 & ~n729;
  assign n731 = ~259 & n729;
  assign n732 = ~n730 & ~n731;
  assign n733 = ~16 & 19;
  assign n734 = 16 & ~n470;
  assign n735 = ~n733 & ~n734;
  assign n736 = 256 & ~n735;
  assign n737 = ~256 & n735;
  assign n738 = ~n736 & ~n737;
  assign n739 = n714 & n720;
  assign n740 = n726 & n739;
  assign n741 = n732 & n740;
  assign n742 = n738 & n741;
  assign n743 = n708 & n742;
  assign n744 = 28 & ~29;
  assign n745 = 29 & ~n567;
  assign n746 = ~n744 & ~n745;
  assign n747 = ~29 & 35;
  assign n748 = 29 & ~1817;
  assign n749 = ~n747 & ~n748;
  assign n750 = 309 & ~n749;
  assign n751 = ~309 & n749;
  assign n752 = ~n750 & ~n751;
  assign n753 = ~n746 & n752;
  assign n754 = ~29 & 34;
  assign n755 = 29 & ~1816;
  assign n756 = ~n754 & ~n755;
  assign n757 = 305 & ~n756;
  assign n758 = ~305 & n756;
  assign n759 = ~n757 & ~n758;
  assign n760 = 27 & ~29;
  assign n761 = 29 & ~1818;
  assign n762 = ~n760 & ~n761;
  assign n763 = 301 & ~n762;
  assign n764 = ~301 & n762;
  assign n765 = ~n763 & ~n764;
  assign n766 = ~29 & 33;
  assign n767 = 139 & ~319;
  assign n768 = ~322 & n767;
  assign n769 = 103 & 319;
  assign n770 = ~322 & n769;
  assign n771 = 127 & ~319;
  assign n772 = 322 & n771;
  assign n773 = 115 & 319;
  assign n774 = 322 & n773;
  assign n775 = ~n768 & ~n770;
  assign n776 = ~n772 & n775;
  assign n777 = ~n774 & n776;
  assign n778 = 29 & ~n777;
  assign n779 = ~n766 & ~n778;
  assign n780 = 297 & ~n779;
  assign n781 = ~297 & n779;
  assign n782 = ~n780 & ~n781;
  assign n783 = 26 & ~29;
  assign n784 = 140 & ~319;
  assign n785 = ~322 & n784;
  assign n786 = 104 & 319;
  assign n787 = ~322 & n786;
  assign n788 = 128 & ~319;
  assign n789 = 322 & n788;
  assign n790 = 116 & 319;
  assign n791 = 322 & n790;
  assign n792 = ~n785 & ~n787;
  assign n793 = ~n789 & n792;
  assign n794 = ~n791 & n793;
  assign n795 = 29 & ~n794;
  assign n796 = ~n783 & ~n795;
  assign n797 = 294 & ~n796;
  assign n798 = ~294 & n796;
  assign n799 = ~n797 & ~n798;
  assign n800 = ~29 & 32;
  assign n801 = 141 & ~319;
  assign n802 = ~322 & n801;
  assign n803 = 105 & 319;
  assign n804 = ~322 & n803;
  assign n805 = 129 & ~319;
  assign n806 = 322 & n805;
  assign n807 = 117 & 319;
  assign n808 = 322 & n807;
  assign n809 = ~n802 & ~n804;
  assign n810 = ~n806 & n809;
  assign n811 = ~n808 & n810;
  assign n812 = 29 & ~n811;
  assign n813 = ~n800 & ~n812;
  assign n814 = 287 & ~n813;
  assign n815 = ~287 & n813;
  assign n816 = ~n814 & ~n815;
  assign n817 = n759 & n765;
  assign n818 = n782 & n817;
  assign n819 = n799 & n818;
  assign n820 = n816 & n819;
  assign n821 = n753 & n820;
  assign n822 = 11 & ~246;
  assign n823 = 11 & 246;
  assign n824 = ~n822 & ~n823;
  assign n825 = n743 & n821;
  assign 3038 = ~n824 & n825;
  assign n827 = ~n470 & n532;
  assign n828 = n470 & ~n532;
  assign n829 = ~n827 & ~n828;
  assign n830 = ~n539 & ~n829;
  assign n831 = n539 & n829;
  assign n832 = ~n830 & ~n831;
  assign n833 = 93 & ~227;
  assign n834 = ~234 & n833;
  assign n835 = 55 & 227;
  assign n836 = ~234 & n835;
  assign n837 = 67 & ~227;
  assign n838 = 234 & n837;
  assign n839 = 80 & 227;
  assign n840 = 234 & n839;
  assign n841 = ~n834 & ~n836;
  assign n842 = ~n838 & n841;
  assign n843 = ~n840 & n842;
  assign n844 = ~n832 & n843;
  assign n845 = n832 & ~n843;
  assign n846 = ~n844 & ~n845;
  assign n847 = ~241 & ~n846;
  assign n848 = 241 & ~n843;
  assign 3546 = n847 | n848;
  assign n850 = ~1816 & 1817;
  assign n851 = 1816 & ~1817;
  assign n852 = ~n850 & ~n851;
  assign n853 = n552 & ~n567;
  assign n854 = ~n552 & n567;
  assign n855 = ~n853 & ~n854;
  assign n856 = ~n852 & n855;
  assign n857 = n852 & ~n855;
  assign n858 = ~n856 & ~n857;
  assign n859 = 142 & ~319;
  assign n860 = ~322 & n859;
  assign n861 = 106 & 319;
  assign n862 = ~322 & n861;
  assign n863 = 130 & ~319;
  assign n864 = 322 & n863;
  assign n865 = 118 & 319;
  assign n866 = 322 & n865;
  assign n867 = ~n860 & ~n862;
  assign n868 = ~n864 & n867;
  assign n869 = ~n866 & n868;
  assign n870 = n675 & ~n869;
  assign n871 = ~n675 & n869;
  assign n872 = ~n870 & ~n871;
  assign n873 = n794 & ~n811;
  assign n874 = ~n794 & n811;
  assign n875 = ~n873 & ~n874;
  assign n876 = 1818 & ~n777;
  assign n877 = ~1818 & n777;
  assign n878 = ~n876 & ~n877;
  assign n879 = ~n872 & n875;
  assign n880 = n878 & n879;
  assign n881 = n872 & n875;
  assign n882 = ~n878 & n881;
  assign n883 = ~n880 & ~n882;
  assign n884 = n872 & ~n875;
  assign n885 = n878 & n884;
  assign n886 = ~n872 & ~n875;
  assign n887 = ~n878 & n886;
  assign n888 = ~n885 & ~n887;
  assign n889 = n883 & n888;
  assign n890 = ~n858 & n889;
  assign n891 = n858 & ~n889;
  assign n892 = ~n890 & ~n891;
  assign 3671 = ~37 & n892;
  assign n894 = ~246 & ~n843;
  assign n895 = 1819 & 2018;
  assign n896 = ~1819 & ~2018;
  assign n897 = ~n895 & ~n896;
  assign n898 = ~2020 & 2022;
  assign n899 = 2020 & ~2022;
  assign n900 = ~n898 & ~n899;
  assign n901 = ~n897 & n900;
  assign n902 = n897 & ~n900;
  assign n903 = ~n901 & ~n902;
  assign n904 = ~n470 & n843;
  assign n905 = n470 & ~n843;
  assign n906 = ~n904 & ~n905;
  assign n907 = 2010 & n532;
  assign n908 = ~2010 & ~n532;
  assign n909 = ~n907 & ~n908;
  assign n910 = ~n539 & n906;
  assign n911 = n909 & n910;
  assign n912 = n539 & n906;
  assign n913 = ~n909 & n912;
  assign n914 = ~n911 & ~n913;
  assign n915 = n539 & ~n906;
  assign n916 = n909 & n915;
  assign n917 = ~n539 & ~n906;
  assign n918 = ~n909 & n917;
  assign n919 = ~n916 & ~n918;
  assign n920 = n914 & n919;
  assign n921 = ~n903 & n920;
  assign n922 = n903 & ~n920;
  assign n923 = ~n921 & ~n922;
  assign n924 = 246 & ~n923;
  assign 3803 = n894 | n924;
  assign n926 = ~1820 & 1821;
  assign n927 = 1820 & ~1821;
  assign n928 = ~n926 & ~n927;
  assign n929 = ~n906 & n909;
  assign n930 = n928 & n929;
  assign n931 = n906 & n909;
  assign n932 = ~n928 & n931;
  assign n933 = ~n930 & ~n932;
  assign n934 = n906 & ~n909;
  assign n935 = n928 & n934;
  assign n936 = ~n906 & ~n909;
  assign n937 = ~n928 & n936;
  assign n938 = ~n935 & ~n937;
  assign n939 = n933 & n938;
  assign n940 = ~n903 & n939;
  assign n941 = n903 & ~n939;
  assign n942 = ~n940 & ~n941;
  assign 3809 = ~37 & n942;
  assign n944 = ~262 & ~1818;
  assign n945 = 1816 & n944;
  assign n946 = 40 & n945;
  assign n947 = ~294 & ~n946;
  assign n948 = 40 & 1816;
  assign n949 = ~n944 & n948;
  assign n950 = n947 & n949;
  assign n951 = ~n794 & ~n946;
  assign n952 = n949 & n951;
  assign n953 = n950 & ~n952;
  assign n954 = ~n950 & ~n952;
  assign n955 = n950 & n952;
  assign n956 = ~n954 & ~n955;
  assign n957 = ~287 & ~n946;
  assign n958 = n949 & n957;
  assign n959 = ~n811 & ~n946;
  assign n960 = n949 & n959;
  assign n961 = n958 & ~n960;
  assign n962 = ~n956 & n961;
  assign n963 = ~n958 & ~n960;
  assign n964 = n958 & n960;
  assign n965 = ~n963 & ~n964;
  assign n966 = ~284 & ~n946;
  assign n967 = n949 & n966;
  assign n968 = ~n675 & ~n946;
  assign n969 = n949 & n968;
  assign n970 = n967 & ~n969;
  assign n971 = ~n956 & ~n965;
  assign n972 = n970 & n971;
  assign n973 = ~n967 & ~n969;
  assign n974 = n967 & n969;
  assign n975 = ~n973 & ~n974;
  assign n976 = 2022 & ~n946;
  assign n977 = n949 & n976;
  assign n978 = ~281 & ~n946;
  assign n979 = n949 & n978;
  assign n980 = ~n977 & n979;
  assign n981 = ~n956 & ~n975;
  assign n982 = n980 & n981;
  assign n983 = ~n965 & n982;
  assign n984 = ~n953 & ~n962;
  assign n985 = ~n972 & n984;
  assign n986 = ~n983 & n985;
  assign n987 = ~278 & ~n946;
  assign n988 = 8 & n987;
  assign n989 = 2020 & ~n946;
  assign n990 = 8 & n989;
  assign n991 = n988 & ~n990;
  assign n992 = ~n988 & ~n990;
  assign n993 = n988 & n990;
  assign n994 = ~n992 & ~n993;
  assign n995 = ~275 & ~n946;
  assign n996 = 8 & n995;
  assign n997 = 2018 & ~n946;
  assign n998 = 8 & n997;
  assign n999 = n996 & ~n998;
  assign n1000 = ~n994 & n999;
  assign n1001 = ~n996 & ~n998;
  assign n1002 = n996 & n998;
  assign n1003 = ~n1001 & ~n1002;
  assign n1004 = ~309 & n946;
  assign n1005 = ~272 & ~n946;
  assign n1006 = ~n1004 & ~n1005;
  assign n1007 = 8 & ~n1006;
  assign n1008 = ~1819 & ~n946;
  assign n1009 = ~1819 & n946;
  assign n1010 = ~n1008 & ~n1009;
  assign n1011 = 8 & ~n1010;
  assign n1012 = n1007 & ~n1011;
  assign n1013 = ~n994 & ~n1003;
  assign n1014 = n1012 & n1013;
  assign n1015 = ~n1007 & ~n1011;
  assign n1016 = n1007 & n1011;
  assign n1017 = ~n1015 & ~n1016;
  assign n1018 = ~305 & n946;
  assign n1019 = ~269 & ~n946;
  assign n1020 = ~n1018 & ~n1019;
  assign n1021 = 8 & ~n1020;
  assign n1022 = ~1820 & ~n946;
  assign n1023 = ~1820 & n946;
  assign n1024 = ~n1022 & ~n1023;
  assign n1025 = 8 & ~n1024;
  assign n1026 = n1021 & ~n1025;
  assign n1027 = ~n994 & ~n1017;
  assign n1028 = n1026 & n1027;
  assign n1029 = ~n1003 & n1028;
  assign n1030 = ~n1021 & ~n1025;
  assign n1031 = n1021 & n1025;
  assign n1032 = ~n1030 & ~n1031;
  assign n1033 = ~301 & n946;
  assign n1034 = ~266 & ~n946;
  assign n1035 = ~n1033 & ~n1034;
  assign n1036 = 1821 & ~n1035;
  assign n1037 = ~n1017 & ~n1032;
  assign n1038 = ~n994 & n1037;
  assign n1039 = n1036 & n1038;
  assign n1040 = ~n1003 & n1039;
  assign n1041 = ~n991 & ~n1000;
  assign n1042 = ~n1014 & n1041;
  assign n1043 = ~n1029 & n1042;
  assign n1044 = ~n1040 & n1043;
  assign n1045 = 1821 & n1035;
  assign n1046 = ~1821 & ~n1035;
  assign n1047 = ~n1045 & ~n1046;
  assign n1048 = ~n1003 & ~n1047;
  assign n1049 = ~n1017 & n1048;
  assign n1050 = ~n994 & n1049;
  assign n1051 = ~n1032 & n1050;
  assign n1052 = ~297 & n946;
  assign n1053 = ~263 & ~n946;
  assign n1054 = ~n1052 & ~n1053;
  assign n1055 = ~2010 & ~n1054;
  assign n1056 = ~2010 & n1054;
  assign n1057 = 2010 & ~n1054;
  assign n1058 = ~n1056 & ~n1057;
  assign n1059 = ~294 & n946;
  assign n1060 = ~259 & ~n946;
  assign n1061 = ~n1059 & ~n1060;
  assign n1062 = n532 & ~n1061;
  assign n1063 = ~n1058 & n1062;
  assign n1064 = n532 & n1061;
  assign n1065 = ~n532 & ~n1061;
  assign n1066 = ~n1064 & ~n1065;
  assign n1067 = ~287 & n946;
  assign n1068 = ~256 & ~n946;
  assign n1069 = ~n1067 & ~n1068;
  assign n1070 = n470 & ~n1069;
  assign n1071 = ~n1058 & ~n1066;
  assign n1072 = n1070 & n1071;
  assign n1073 = ~n1055 & ~n1063;
  assign n1074 = ~n1072 & n1073;
  assign n1075 = n1051 & ~n1074;
  assign n1076 = n1044 & ~n1075;
  assign n1077 = ~n986 & n1076;
  assign n1078 = ~n977 & ~n979;
  assign n1079 = n977 & n979;
  assign n1080 = ~n1078 & ~n1079;
  assign n1081 = ~n965 & ~n1080;
  assign n1082 = ~n975 & n1081;
  assign n1083 = ~n956 & n1082;
  assign n1084 = n986 & ~n1083;
  assign n1085 = ~n1076 & ~n1084;
  assign 3851 = n1077 | n1085;
  assign n1087 = ~3671 & ~3809;
  assign n1088 = ~2970 & n1087;
  assign n1089 = ~2925 & ~2971;
  assign n1090 = n1088 & n1089;
  assign 3881 = 1726 & n1090;
  assign 3875 = 1'b0;
  assign 487 = ~44;
  assign 488 = ~132;
  assign 489 = ~82;
  assign 490 = ~96;
  assign 491 = ~69;
  assign 492 = ~120;
  assign 493 = ~57;
  assign 494 = ~108;
  assign 1448 = ~1277;
  assign 2012 = ~1821;
  assign 2014 = ~1820;
  assign 2016 = ~1819;
  assign 3079 = ~3038;
  assign 3882 = ~3881;
  assign 398 = 219;
  assign 400 = 219;
  assign 401 = 219;
  assign 419 = 253;
  assign 420 = 253;
  assign 456 = 290;
  assign 457 = 290;
  assign 458 = 290;
  assign 805 = 219;
  assign 2388 = 2387;
  assign 2390 = 2389;
  assign 2644 = 2643;
  assign 3804 = 3803;
endmodule
