module top (
    \1 , 18, 35, 52, 69, 86, 103, 120, 137, 154, 171, 188, 205, 222, 239,
    256, 273, 290, 307, 324, 341, 358, 375, 392, 409, 426, 443, 460, 477,
    494, 511, 528,
    545, 1581, 1901, 2223, 2548, 2877, 3211, 3552, 3895, 4241, 4591, 4946,
    5308, 5672, 5971, 6123, 6150, 6160, 6170, 6180, 6190, 6200, 6210, 6220,
    6230, 6240, 6250, 6260, 6270, 6280, 6287, 6288  );
  input  \1 , 18, 35, 52, 69, 86, 103, 120, 137, 154, 171, 188, 205, 222,
    239, 256, 273, 290, 307, 324, 341, 358, 375, 392, 409, 426, 443, 460,
    477, 494, 511, 528;
  output 545, 1581, 1901, 2223, 2548, 2877, 3211, 3552, 3895, 4241, 4591,
    4946, 5308, 5672, 5971, 6123, 6150, 6160, 6170, 6180, 6190, 6200, 6210,
    6220, 6230, 6240, 6250, 6260, 6270, 6280, 6287, 6288;
  wire n66, n67, n68, n69, n70, n72, n73, n74, n75, n76, n77, n78, n79, n80,
    n81, n82, n83, n84, n85, n87, n88, n89, n90, n91, n92, n93, n94, n95,
    n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107,
    n108, n109, n110, n112, n113, n114, n115, n116, n117, n118, n119, n120,
    n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
    n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
    n145, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157,
    n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169,
    n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181,
    n182, n183, n184, n185, n186, n187, n188, n189, n190, n192, n193, n194,
    n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206,
    n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218,
    n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230,
    n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
    n243, n244, n245, n247, n248, n249, n250, n251, n252, n253, n254, n255,
    n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267,
    n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
    n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291,
    n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
    n304, n305, n306, n307, n308, n309, n310, n312, n313, n314, n315, n316,
    n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328,
    n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340,
    n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
    n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
    n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
    n377, n378, n379, n380, n381, n382, n383, n384, n385, n387, n388, n389,
    n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
    n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
    n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
    n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
    n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
    n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
    n462, n463, n464, n465, n466, n467, n468, n469, n470, n472, n473, n474,
    n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
    n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
    n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
    n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
    n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
    n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
    n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
    n559, n560, n561, n562, n563, n564, n565, n567, n568, n569, n570, n571,
    n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
    n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
    n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
    n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
    n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
    n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
    n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
    n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
    n668, n669, n670, n672, n673, n674, n675, n676, n677, n678, n679, n680,
    n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
    n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
    n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
    n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
    n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
    n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
    n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764,
    n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
    n777, n778, n779, n780, n781, n782, n783, n784, n785, n787, n788, n789,
    n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
    n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813,
    n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825,
    n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
    n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
    n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
    n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873,
    n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885,
    n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897,
    n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909,
    n910, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922,
    n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934,
    n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946,
    n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
    n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
    n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
    n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
    n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005,
    n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
    n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
    n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035,
    n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045,
    n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056,
    n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066,
    n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076,
    n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086,
    n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096,
    n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106,
    n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116,
    n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126,
    n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136,
    n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146,
    n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156,
    n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166,
    n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176,
    n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186,
    n1187, n1188, n1189, n1190, n1192, n1193, n1194, n1195, n1196, n1197,
    n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207,
    n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217,
    n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227,
    n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237,
    n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247,
    n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257,
    n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267,
    n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277,
    n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287,
    n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297,
    n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307,
    n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317,
    n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327,
    n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1337, n1338,
    n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348,
    n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358,
    n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368,
    n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378,
    n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388,
    n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398,
    n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408,
    n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418,
    n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428,
    n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438,
    n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448,
    n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458,
    n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468,
    n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1478, n1479,
    n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489,
    n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499,
    n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509,
    n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519,
    n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529,
    n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539,
    n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549,
    n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559,
    n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569,
    n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579,
    n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589,
    n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599,
    n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1609, n1610,
    n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620,
    n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630,
    n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640,
    n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650,
    n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660,
    n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670,
    n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680,
    n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690,
    n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700,
    n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710,
    n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720,
    n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1730, n1731,
    n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741,
    n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751,
    n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761,
    n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771,
    n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781,
    n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791,
    n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801,
    n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811,
    n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821,
    n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831,
    n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1841, n1842,
    n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
    n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
    n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
    n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
    n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
    n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
    n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
    n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
    n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
    n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1942, n1943,
    n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953,
    n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963,
    n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973,
    n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983,
    n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993,
    n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003,
    n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013,
    n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023,
    n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2033, n2034,
    n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044,
    n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054,
    n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064,
    n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074,
    n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084,
    n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094,
    n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104,
    n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2114, n2115,
    n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125,
    n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135,
    n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145,
    n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155,
    n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165,
    n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175,
    n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2185, n2186,
    n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196,
    n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206,
    n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216,
    n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226,
    n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236,
    n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2246, n2247,
    n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257,
    n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267,
    n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277,
    n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287,
    n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2297, n2298,
    n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308,
    n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318,
    n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328,
    n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2338, n2339,
    n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349,
    n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359,
    n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2369, n2370,
    n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380,
    n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2390, n2391,
    n2392, n2393, n2394, n2395, n2396, n2397, n2399, n2400;
  assign 545 = \1  & 273;
  assign n66 = 18 & 273;
  assign n67 = \1  & 290;
  assign n68 = n66 & ~n67;
  assign n69 = n66 & ~n68;
  assign n70 = ~n67 & ~n68;
  assign 1581 = ~n69 & ~n70;
  assign n72 = 35 & 273;
  assign n73 = 18 & 290;
  assign n74 = n72 & ~n73;
  assign n75 = n72 & ~n74;
  assign n76 = ~n73 & ~n74;
  assign n77 = ~n75 & ~n76;
  assign n78 = ~n69 & ~n77;
  assign n79 = ~n77 & ~n78;
  assign n80 = ~n69 & ~n78;
  assign n81 = ~n79 & ~n80;
  assign n82 = \1  & 307;
  assign n83 = ~n81 & ~n82;
  assign n84 = ~n81 & ~n83;
  assign n85 = ~n82 & ~n83;
  assign 1901 = ~n84 & ~n85;
  assign n87 = 52 & 273;
  assign n88 = 35 & 290;
  assign n89 = n87 & ~n88;
  assign n90 = n87 & ~n89;
  assign n91 = ~n88 & ~n89;
  assign n92 = ~n90 & ~n91;
  assign n93 = ~n75 & ~n92;
  assign n94 = ~n92 & ~n93;
  assign n95 = ~n75 & ~n93;
  assign n96 = ~n94 & ~n95;
  assign n97 = 18 & 307;
  assign n98 = ~n96 & ~n97;
  assign n99 = ~n96 & ~n98;
  assign n100 = ~n97 & ~n98;
  assign n101 = ~n99 & ~n100;
  assign n102 = ~n78 & ~n83;
  assign n103 = ~n101 & ~n102;
  assign n104 = ~n101 & ~n103;
  assign n105 = ~n102 & ~n103;
  assign n106 = ~n104 & ~n105;
  assign n107 = \1  & 324;
  assign n108 = ~n106 & ~n107;
  assign n109 = ~n106 & ~n108;
  assign n110 = ~n107 & ~n108;
  assign 2223 = ~n109 & ~n110;
  assign n112 = 69 & 273;
  assign n113 = 52 & 290;
  assign n114 = n112 & ~n113;
  assign n115 = n112 & ~n114;
  assign n116 = ~n113 & ~n114;
  assign n117 = ~n115 & ~n116;
  assign n118 = ~n90 & ~n117;
  assign n119 = ~n117 & ~n118;
  assign n120 = ~n90 & ~n118;
  assign n121 = ~n119 & ~n120;
  assign n122 = 35 & 307;
  assign n123 = ~n121 & ~n122;
  assign n124 = ~n121 & ~n123;
  assign n125 = ~n122 & ~n123;
  assign n126 = ~n124 & ~n125;
  assign n127 = ~n93 & ~n98;
  assign n128 = ~n126 & ~n127;
  assign n129 = ~n126 & ~n128;
  assign n130 = ~n127 & ~n128;
  assign n131 = ~n129 & ~n130;
  assign n132 = 18 & 324;
  assign n133 = ~n131 & ~n132;
  assign n134 = ~n131 & ~n133;
  assign n135 = ~n132 & ~n133;
  assign n136 = ~n134 & ~n135;
  assign n137 = ~n103 & ~n108;
  assign n138 = ~n136 & ~n137;
  assign n139 = ~n136 & ~n138;
  assign n140 = ~n137 & ~n138;
  assign n141 = ~n139 & ~n140;
  assign n142 = \1  & 341;
  assign n143 = ~n141 & ~n142;
  assign n144 = ~n141 & ~n143;
  assign n145 = ~n142 & ~n143;
  assign 2548 = ~n144 & ~n145;
  assign n147 = 86 & 273;
  assign n148 = 69 & 290;
  assign n149 = n147 & ~n148;
  assign n150 = n147 & ~n149;
  assign n151 = ~n148 & ~n149;
  assign n152 = ~n150 & ~n151;
  assign n153 = ~n115 & ~n152;
  assign n154 = ~n152 & ~n153;
  assign n155 = ~n115 & ~n153;
  assign n156 = ~n154 & ~n155;
  assign n157 = 52 & 307;
  assign n158 = ~n156 & ~n157;
  assign n159 = ~n156 & ~n158;
  assign n160 = ~n157 & ~n158;
  assign n161 = ~n159 & ~n160;
  assign n162 = ~n118 & ~n123;
  assign n163 = ~n161 & ~n162;
  assign n164 = ~n161 & ~n163;
  assign n165 = ~n162 & ~n163;
  assign n166 = ~n164 & ~n165;
  assign n167 = 35 & 324;
  assign n168 = ~n166 & ~n167;
  assign n169 = ~n166 & ~n168;
  assign n170 = ~n167 & ~n168;
  assign n171 = ~n169 & ~n170;
  assign n172 = ~n128 & ~n133;
  assign n173 = ~n171 & ~n172;
  assign n174 = ~n171 & ~n173;
  assign n175 = ~n172 & ~n173;
  assign n176 = ~n174 & ~n175;
  assign n177 = 18 & 341;
  assign n178 = ~n176 & ~n177;
  assign n179 = ~n176 & ~n178;
  assign n180 = ~n177 & ~n178;
  assign n181 = ~n179 & ~n180;
  assign n182 = ~n138 & ~n143;
  assign n183 = ~n181 & ~n182;
  assign n184 = ~n181 & ~n183;
  assign n185 = ~n182 & ~n183;
  assign n186 = ~n184 & ~n185;
  assign n187 = \1  & 358;
  assign n188 = ~n186 & ~n187;
  assign n189 = ~n186 & ~n188;
  assign n190 = ~n187 & ~n188;
  assign 2877 = ~n189 & ~n190;
  assign n192 = 103 & 273;
  assign n193 = 86 & 290;
  assign n194 = n192 & ~n193;
  assign n195 = n192 & ~n194;
  assign n196 = ~n193 & ~n194;
  assign n197 = ~n195 & ~n196;
  assign n198 = ~n150 & ~n197;
  assign n199 = ~n197 & ~n198;
  assign n200 = ~n150 & ~n198;
  assign n201 = ~n199 & ~n200;
  assign n202 = 69 & 307;
  assign n203 = ~n201 & ~n202;
  assign n204 = ~n201 & ~n203;
  assign n205 = ~n202 & ~n203;
  assign n206 = ~n204 & ~n205;
  assign n207 = ~n153 & ~n158;
  assign n208 = ~n206 & ~n207;
  assign n209 = ~n206 & ~n208;
  assign n210 = ~n207 & ~n208;
  assign n211 = ~n209 & ~n210;
  assign n212 = 52 & 324;
  assign n213 = ~n211 & ~n212;
  assign n214 = ~n211 & ~n213;
  assign n215 = ~n212 & ~n213;
  assign n216 = ~n214 & ~n215;
  assign n217 = ~n163 & ~n168;
  assign n218 = ~n216 & ~n217;
  assign n219 = ~n216 & ~n218;
  assign n220 = ~n217 & ~n218;
  assign n221 = ~n219 & ~n220;
  assign n222 = 35 & 341;
  assign n223 = ~n221 & ~n222;
  assign n224 = ~n221 & ~n223;
  assign n225 = ~n222 & ~n223;
  assign n226 = ~n224 & ~n225;
  assign n227 = ~n173 & ~n178;
  assign n228 = ~n226 & ~n227;
  assign n229 = ~n226 & ~n228;
  assign n230 = ~n227 & ~n228;
  assign n231 = ~n229 & ~n230;
  assign n232 = 18 & 358;
  assign n233 = ~n231 & ~n232;
  assign n234 = ~n231 & ~n233;
  assign n235 = ~n232 & ~n233;
  assign n236 = ~n234 & ~n235;
  assign n237 = ~n183 & ~n188;
  assign n238 = ~n236 & ~n237;
  assign n239 = ~n236 & ~n238;
  assign n240 = ~n237 & ~n238;
  assign n241 = ~n239 & ~n240;
  assign n242 = \1  & 375;
  assign n243 = ~n241 & ~n242;
  assign n244 = ~n241 & ~n243;
  assign n245 = ~n242 & ~n243;
  assign 3211 = ~n244 & ~n245;
  assign n247 = 120 & 273;
  assign n248 = 103 & 290;
  assign n249 = n247 & ~n248;
  assign n250 = n247 & ~n249;
  assign n251 = ~n248 & ~n249;
  assign n252 = ~n250 & ~n251;
  assign n253 = ~n195 & ~n252;
  assign n254 = ~n252 & ~n253;
  assign n255 = ~n195 & ~n253;
  assign n256 = ~n254 & ~n255;
  assign n257 = 86 & 307;
  assign n258 = ~n256 & ~n257;
  assign n259 = ~n256 & ~n258;
  assign n260 = ~n257 & ~n258;
  assign n261 = ~n259 & ~n260;
  assign n262 = ~n198 & ~n203;
  assign n263 = ~n261 & ~n262;
  assign n264 = ~n261 & ~n263;
  assign n265 = ~n262 & ~n263;
  assign n266 = ~n264 & ~n265;
  assign n267 = 69 & 324;
  assign n268 = ~n266 & ~n267;
  assign n269 = ~n266 & ~n268;
  assign n270 = ~n267 & ~n268;
  assign n271 = ~n269 & ~n270;
  assign n272 = ~n208 & ~n213;
  assign n273 = ~n271 & ~n272;
  assign n274 = ~n271 & ~n273;
  assign n275 = ~n272 & ~n273;
  assign n276 = ~n274 & ~n275;
  assign n277 = 52 & 341;
  assign n278 = ~n276 & ~n277;
  assign n279 = ~n276 & ~n278;
  assign n280 = ~n277 & ~n278;
  assign n281 = ~n279 & ~n280;
  assign n282 = ~n218 & ~n223;
  assign n283 = ~n281 & ~n282;
  assign n284 = ~n281 & ~n283;
  assign n285 = ~n282 & ~n283;
  assign n286 = ~n284 & ~n285;
  assign n287 = 35 & 358;
  assign n288 = ~n286 & ~n287;
  assign n289 = ~n286 & ~n288;
  assign n290 = ~n287 & ~n288;
  assign n291 = ~n289 & ~n290;
  assign n292 = ~n228 & ~n233;
  assign n293 = ~n291 & ~n292;
  assign n294 = ~n291 & ~n293;
  assign n295 = ~n292 & ~n293;
  assign n296 = ~n294 & ~n295;
  assign n297 = 18 & 375;
  assign n298 = ~n296 & ~n297;
  assign n299 = ~n296 & ~n298;
  assign n300 = ~n297 & ~n298;
  assign n301 = ~n299 & ~n300;
  assign n302 = ~n238 & ~n243;
  assign n303 = ~n301 & ~n302;
  assign n304 = ~n301 & ~n303;
  assign n305 = ~n302 & ~n303;
  assign n306 = ~n304 & ~n305;
  assign n307 = \1  & 392;
  assign n308 = ~n306 & ~n307;
  assign n309 = ~n306 & ~n308;
  assign n310 = ~n307 & ~n308;
  assign 3552 = ~n309 & ~n310;
  assign n312 = 137 & 273;
  assign n313 = 120 & 290;
  assign n314 = n312 & ~n313;
  assign n315 = n312 & ~n314;
  assign n316 = ~n313 & ~n314;
  assign n317 = ~n315 & ~n316;
  assign n318 = ~n250 & ~n317;
  assign n319 = ~n317 & ~n318;
  assign n320 = ~n250 & ~n318;
  assign n321 = ~n319 & ~n320;
  assign n322 = 103 & 307;
  assign n323 = ~n321 & ~n322;
  assign n324 = ~n321 & ~n323;
  assign n325 = ~n322 & ~n323;
  assign n326 = ~n324 & ~n325;
  assign n327 = ~n253 & ~n258;
  assign n328 = ~n326 & ~n327;
  assign n329 = ~n326 & ~n328;
  assign n330 = ~n327 & ~n328;
  assign n331 = ~n329 & ~n330;
  assign n332 = 86 & 324;
  assign n333 = ~n331 & ~n332;
  assign n334 = ~n331 & ~n333;
  assign n335 = ~n332 & ~n333;
  assign n336 = ~n334 & ~n335;
  assign n337 = ~n263 & ~n268;
  assign n338 = ~n336 & ~n337;
  assign n339 = ~n336 & ~n338;
  assign n340 = ~n337 & ~n338;
  assign n341 = ~n339 & ~n340;
  assign n342 = 69 & 341;
  assign n343 = ~n341 & ~n342;
  assign n344 = ~n341 & ~n343;
  assign n345 = ~n342 & ~n343;
  assign n346 = ~n344 & ~n345;
  assign n347 = ~n273 & ~n278;
  assign n348 = ~n346 & ~n347;
  assign n349 = ~n346 & ~n348;
  assign n350 = ~n347 & ~n348;
  assign n351 = ~n349 & ~n350;
  assign n352 = 52 & 358;
  assign n353 = ~n351 & ~n352;
  assign n354 = ~n351 & ~n353;
  assign n355 = ~n352 & ~n353;
  assign n356 = ~n354 & ~n355;
  assign n357 = ~n283 & ~n288;
  assign n358 = ~n356 & ~n357;
  assign n359 = ~n356 & ~n358;
  assign n360 = ~n357 & ~n358;
  assign n361 = ~n359 & ~n360;
  assign n362 = 35 & 375;
  assign n363 = ~n361 & ~n362;
  assign n364 = ~n361 & ~n363;
  assign n365 = ~n362 & ~n363;
  assign n366 = ~n364 & ~n365;
  assign n367 = ~n293 & ~n298;
  assign n368 = ~n366 & ~n367;
  assign n369 = ~n366 & ~n368;
  assign n370 = ~n367 & ~n368;
  assign n371 = ~n369 & ~n370;
  assign n372 = 18 & 392;
  assign n373 = ~n371 & ~n372;
  assign n374 = ~n371 & ~n373;
  assign n375 = ~n372 & ~n373;
  assign n376 = ~n374 & ~n375;
  assign n377 = ~n303 & ~n308;
  assign n378 = ~n376 & ~n377;
  assign n379 = ~n376 & ~n378;
  assign n380 = ~n377 & ~n378;
  assign n381 = ~n379 & ~n380;
  assign n382 = \1  & 409;
  assign n383 = ~n381 & ~n382;
  assign n384 = ~n381 & ~n383;
  assign n385 = ~n382 & ~n383;
  assign 3895 = ~n384 & ~n385;
  assign n387 = 154 & 273;
  assign n388 = 137 & 290;
  assign n389 = n387 & ~n388;
  assign n390 = n387 & ~n389;
  assign n391 = ~n388 & ~n389;
  assign n392 = ~n390 & ~n391;
  assign n393 = ~n315 & ~n392;
  assign n394 = ~n392 & ~n393;
  assign n395 = ~n315 & ~n393;
  assign n396 = ~n394 & ~n395;
  assign n397 = 120 & 307;
  assign n398 = ~n396 & ~n397;
  assign n399 = ~n396 & ~n398;
  assign n400 = ~n397 & ~n398;
  assign n401 = ~n399 & ~n400;
  assign n402 = ~n318 & ~n323;
  assign n403 = ~n401 & ~n402;
  assign n404 = ~n401 & ~n403;
  assign n405 = ~n402 & ~n403;
  assign n406 = ~n404 & ~n405;
  assign n407 = 103 & 324;
  assign n408 = ~n406 & ~n407;
  assign n409 = ~n406 & ~n408;
  assign n410 = ~n407 & ~n408;
  assign n411 = ~n409 & ~n410;
  assign n412 = ~n328 & ~n333;
  assign n413 = ~n411 & ~n412;
  assign n414 = ~n411 & ~n413;
  assign n415 = ~n412 & ~n413;
  assign n416 = ~n414 & ~n415;
  assign n417 = 86 & 341;
  assign n418 = ~n416 & ~n417;
  assign n419 = ~n416 & ~n418;
  assign n420 = ~n417 & ~n418;
  assign n421 = ~n419 & ~n420;
  assign n422 = ~n338 & ~n343;
  assign n423 = ~n421 & ~n422;
  assign n424 = ~n421 & ~n423;
  assign n425 = ~n422 & ~n423;
  assign n426 = ~n424 & ~n425;
  assign n427 = 69 & 358;
  assign n428 = ~n426 & ~n427;
  assign n429 = ~n426 & ~n428;
  assign n430 = ~n427 & ~n428;
  assign n431 = ~n429 & ~n430;
  assign n432 = ~n348 & ~n353;
  assign n433 = ~n431 & ~n432;
  assign n434 = ~n431 & ~n433;
  assign n435 = ~n432 & ~n433;
  assign n436 = ~n434 & ~n435;
  assign n437 = 52 & 375;
  assign n438 = ~n436 & ~n437;
  assign n439 = ~n436 & ~n438;
  assign n440 = ~n437 & ~n438;
  assign n441 = ~n439 & ~n440;
  assign n442 = ~n358 & ~n363;
  assign n443 = ~n441 & ~n442;
  assign n444 = ~n441 & ~n443;
  assign n445 = ~n442 & ~n443;
  assign n446 = ~n444 & ~n445;
  assign n447 = 35 & 392;
  assign n448 = ~n446 & ~n447;
  assign n449 = ~n446 & ~n448;
  assign n450 = ~n447 & ~n448;
  assign n451 = ~n449 & ~n450;
  assign n452 = ~n368 & ~n373;
  assign n453 = ~n451 & ~n452;
  assign n454 = ~n451 & ~n453;
  assign n455 = ~n452 & ~n453;
  assign n456 = ~n454 & ~n455;
  assign n457 = 18 & 409;
  assign n458 = ~n456 & ~n457;
  assign n459 = ~n456 & ~n458;
  assign n460 = ~n457 & ~n458;
  assign n461 = ~n459 & ~n460;
  assign n462 = ~n378 & ~n383;
  assign n463 = ~n461 & ~n462;
  assign n464 = ~n461 & ~n463;
  assign n465 = ~n462 & ~n463;
  assign n466 = ~n464 & ~n465;
  assign n467 = \1  & 426;
  assign n468 = ~n466 & ~n467;
  assign n469 = ~n466 & ~n468;
  assign n470 = ~n467 & ~n468;
  assign 4241 = ~n469 & ~n470;
  assign n472 = 171 & 273;
  assign n473 = 154 & 290;
  assign n474 = n472 & ~n473;
  assign n475 = n472 & ~n474;
  assign n476 = ~n473 & ~n474;
  assign n477 = ~n475 & ~n476;
  assign n478 = ~n390 & ~n477;
  assign n479 = ~n477 & ~n478;
  assign n480 = ~n390 & ~n478;
  assign n481 = ~n479 & ~n480;
  assign n482 = 137 & 307;
  assign n483 = ~n481 & ~n482;
  assign n484 = ~n481 & ~n483;
  assign n485 = ~n482 & ~n483;
  assign n486 = ~n484 & ~n485;
  assign n487 = ~n393 & ~n398;
  assign n488 = ~n486 & ~n487;
  assign n489 = ~n486 & ~n488;
  assign n490 = ~n487 & ~n488;
  assign n491 = ~n489 & ~n490;
  assign n492 = 120 & 324;
  assign n493 = ~n491 & ~n492;
  assign n494 = ~n491 & ~n493;
  assign n495 = ~n492 & ~n493;
  assign n496 = ~n494 & ~n495;
  assign n497 = ~n403 & ~n408;
  assign n498 = ~n496 & ~n497;
  assign n499 = ~n496 & ~n498;
  assign n500 = ~n497 & ~n498;
  assign n501 = ~n499 & ~n500;
  assign n502 = 103 & 341;
  assign n503 = ~n501 & ~n502;
  assign n504 = ~n501 & ~n503;
  assign n505 = ~n502 & ~n503;
  assign n506 = ~n504 & ~n505;
  assign n507 = ~n413 & ~n418;
  assign n508 = ~n506 & ~n507;
  assign n509 = ~n506 & ~n508;
  assign n510 = ~n507 & ~n508;
  assign n511 = ~n509 & ~n510;
  assign n512 = 86 & 358;
  assign n513 = ~n511 & ~n512;
  assign n514 = ~n511 & ~n513;
  assign n515 = ~n512 & ~n513;
  assign n516 = ~n514 & ~n515;
  assign n517 = ~n423 & ~n428;
  assign n518 = ~n516 & ~n517;
  assign n519 = ~n516 & ~n518;
  assign n520 = ~n517 & ~n518;
  assign n521 = ~n519 & ~n520;
  assign n522 = 69 & 375;
  assign n523 = ~n521 & ~n522;
  assign n524 = ~n521 & ~n523;
  assign n525 = ~n522 & ~n523;
  assign n526 = ~n524 & ~n525;
  assign n527 = ~n433 & ~n438;
  assign n528 = ~n526 & ~n527;
  assign n529 = ~n526 & ~n528;
  assign n530 = ~n527 & ~n528;
  assign n531 = ~n529 & ~n530;
  assign n532 = 52 & 392;
  assign n533 = ~n531 & ~n532;
  assign n534 = ~n531 & ~n533;
  assign n535 = ~n532 & ~n533;
  assign n536 = ~n534 & ~n535;
  assign n537 = ~n443 & ~n448;
  assign n538 = ~n536 & ~n537;
  assign n539 = ~n536 & ~n538;
  assign n540 = ~n537 & ~n538;
  assign n541 = ~n539 & ~n540;
  assign n542 = 35 & 409;
  assign n543 = ~n541 & ~n542;
  assign n544 = ~n541 & ~n543;
  assign n545 = ~n542 & ~n543;
  assign n546 = ~n544 & ~n545;
  assign n547 = ~n453 & ~n458;
  assign n548 = ~n546 & ~n547;
  assign n549 = ~n546 & ~n548;
  assign n550 = ~n547 & ~n548;
  assign n551 = ~n549 & ~n550;
  assign n552 = 18 & 426;
  assign n553 = ~n551 & ~n552;
  assign n554 = ~n551 & ~n553;
  assign n555 = ~n552 & ~n553;
  assign n556 = ~n554 & ~n555;
  assign n557 = ~n463 & ~n468;
  assign n558 = ~n556 & ~n557;
  assign n559 = ~n556 & ~n558;
  assign n560 = ~n557 & ~n558;
  assign n561 = ~n559 & ~n560;
  assign n562 = \1  & 443;
  assign n563 = ~n561 & ~n562;
  assign n564 = ~n561 & ~n563;
  assign n565 = ~n562 & ~n563;
  assign 4591 = ~n564 & ~n565;
  assign n567 = 188 & 273;
  assign n568 = 171 & 290;
  assign n569 = n567 & ~n568;
  assign n570 = n567 & ~n569;
  assign n571 = ~n568 & ~n569;
  assign n572 = ~n570 & ~n571;
  assign n573 = ~n475 & ~n572;
  assign n574 = ~n572 & ~n573;
  assign n575 = ~n475 & ~n573;
  assign n576 = ~n574 & ~n575;
  assign n577 = 154 & 307;
  assign n578 = ~n576 & ~n577;
  assign n579 = ~n576 & ~n578;
  assign n580 = ~n577 & ~n578;
  assign n581 = ~n579 & ~n580;
  assign n582 = ~n478 & ~n483;
  assign n583 = ~n581 & ~n582;
  assign n584 = ~n581 & ~n583;
  assign n585 = ~n582 & ~n583;
  assign n586 = ~n584 & ~n585;
  assign n587 = 137 & 324;
  assign n588 = ~n586 & ~n587;
  assign n589 = ~n586 & ~n588;
  assign n590 = ~n587 & ~n588;
  assign n591 = ~n589 & ~n590;
  assign n592 = ~n488 & ~n493;
  assign n593 = ~n591 & ~n592;
  assign n594 = ~n591 & ~n593;
  assign n595 = ~n592 & ~n593;
  assign n596 = ~n594 & ~n595;
  assign n597 = 120 & 341;
  assign n598 = ~n596 & ~n597;
  assign n599 = ~n596 & ~n598;
  assign n600 = ~n597 & ~n598;
  assign n601 = ~n599 & ~n600;
  assign n602 = ~n498 & ~n503;
  assign n603 = ~n601 & ~n602;
  assign n604 = ~n601 & ~n603;
  assign n605 = ~n602 & ~n603;
  assign n606 = ~n604 & ~n605;
  assign n607 = 103 & 358;
  assign n608 = ~n606 & ~n607;
  assign n609 = ~n606 & ~n608;
  assign n610 = ~n607 & ~n608;
  assign n611 = ~n609 & ~n610;
  assign n612 = ~n508 & ~n513;
  assign n613 = ~n611 & ~n612;
  assign n614 = ~n611 & ~n613;
  assign n615 = ~n612 & ~n613;
  assign n616 = ~n614 & ~n615;
  assign n617 = 86 & 375;
  assign n618 = ~n616 & ~n617;
  assign n619 = ~n616 & ~n618;
  assign n620 = ~n617 & ~n618;
  assign n621 = ~n619 & ~n620;
  assign n622 = ~n518 & ~n523;
  assign n623 = ~n621 & ~n622;
  assign n624 = ~n621 & ~n623;
  assign n625 = ~n622 & ~n623;
  assign n626 = ~n624 & ~n625;
  assign n627 = 69 & 392;
  assign n628 = ~n626 & ~n627;
  assign n629 = ~n626 & ~n628;
  assign n630 = ~n627 & ~n628;
  assign n631 = ~n629 & ~n630;
  assign n632 = ~n528 & ~n533;
  assign n633 = ~n631 & ~n632;
  assign n634 = ~n631 & ~n633;
  assign n635 = ~n632 & ~n633;
  assign n636 = ~n634 & ~n635;
  assign n637 = 52 & 409;
  assign n638 = ~n636 & ~n637;
  assign n639 = ~n636 & ~n638;
  assign n640 = ~n637 & ~n638;
  assign n641 = ~n639 & ~n640;
  assign n642 = ~n538 & ~n543;
  assign n643 = ~n641 & ~n642;
  assign n644 = ~n641 & ~n643;
  assign n645 = ~n642 & ~n643;
  assign n646 = ~n644 & ~n645;
  assign n647 = 35 & 426;
  assign n648 = ~n646 & ~n647;
  assign n649 = ~n646 & ~n648;
  assign n650 = ~n647 & ~n648;
  assign n651 = ~n649 & ~n650;
  assign n652 = ~n548 & ~n553;
  assign n653 = ~n651 & ~n652;
  assign n654 = ~n651 & ~n653;
  assign n655 = ~n652 & ~n653;
  assign n656 = ~n654 & ~n655;
  assign n657 = 18 & 443;
  assign n658 = ~n656 & ~n657;
  assign n659 = ~n656 & ~n658;
  assign n660 = ~n657 & ~n658;
  assign n661 = ~n659 & ~n660;
  assign n662 = ~n558 & ~n563;
  assign n663 = ~n661 & ~n662;
  assign n664 = ~n661 & ~n663;
  assign n665 = ~n662 & ~n663;
  assign n666 = ~n664 & ~n665;
  assign n667 = \1  & 460;
  assign n668 = ~n666 & ~n667;
  assign n669 = ~n666 & ~n668;
  assign n670 = ~n667 & ~n668;
  assign 4946 = ~n669 & ~n670;
  assign n672 = 205 & 273;
  assign n673 = 188 & 290;
  assign n674 = n672 & ~n673;
  assign n675 = n672 & ~n674;
  assign n676 = ~n673 & ~n674;
  assign n677 = ~n675 & ~n676;
  assign n678 = ~n570 & ~n677;
  assign n679 = ~n677 & ~n678;
  assign n680 = ~n570 & ~n678;
  assign n681 = ~n679 & ~n680;
  assign n682 = 171 & 307;
  assign n683 = ~n681 & ~n682;
  assign n684 = ~n681 & ~n683;
  assign n685 = ~n682 & ~n683;
  assign n686 = ~n684 & ~n685;
  assign n687 = ~n573 & ~n578;
  assign n688 = ~n686 & ~n687;
  assign n689 = ~n686 & ~n688;
  assign n690 = ~n687 & ~n688;
  assign n691 = ~n689 & ~n690;
  assign n692 = 154 & 324;
  assign n693 = ~n691 & ~n692;
  assign n694 = ~n691 & ~n693;
  assign n695 = ~n692 & ~n693;
  assign n696 = ~n694 & ~n695;
  assign n697 = ~n583 & ~n588;
  assign n698 = ~n696 & ~n697;
  assign n699 = ~n696 & ~n698;
  assign n700 = ~n697 & ~n698;
  assign n701 = ~n699 & ~n700;
  assign n702 = 137 & 341;
  assign n703 = ~n701 & ~n702;
  assign n704 = ~n701 & ~n703;
  assign n705 = ~n702 & ~n703;
  assign n706 = ~n704 & ~n705;
  assign n707 = ~n593 & ~n598;
  assign n708 = ~n706 & ~n707;
  assign n709 = ~n706 & ~n708;
  assign n710 = ~n707 & ~n708;
  assign n711 = ~n709 & ~n710;
  assign n712 = 120 & 358;
  assign n713 = ~n711 & ~n712;
  assign n714 = ~n711 & ~n713;
  assign n715 = ~n712 & ~n713;
  assign n716 = ~n714 & ~n715;
  assign n717 = ~n603 & ~n608;
  assign n718 = ~n716 & ~n717;
  assign n719 = ~n716 & ~n718;
  assign n720 = ~n717 & ~n718;
  assign n721 = ~n719 & ~n720;
  assign n722 = 103 & 375;
  assign n723 = ~n721 & ~n722;
  assign n724 = ~n721 & ~n723;
  assign n725 = ~n722 & ~n723;
  assign n726 = ~n724 & ~n725;
  assign n727 = ~n613 & ~n618;
  assign n728 = ~n726 & ~n727;
  assign n729 = ~n726 & ~n728;
  assign n730 = ~n727 & ~n728;
  assign n731 = ~n729 & ~n730;
  assign n732 = 86 & 392;
  assign n733 = ~n731 & ~n732;
  assign n734 = ~n731 & ~n733;
  assign n735 = ~n732 & ~n733;
  assign n736 = ~n734 & ~n735;
  assign n737 = ~n623 & ~n628;
  assign n738 = ~n736 & ~n737;
  assign n739 = ~n736 & ~n738;
  assign n740 = ~n737 & ~n738;
  assign n741 = ~n739 & ~n740;
  assign n742 = 69 & 409;
  assign n743 = ~n741 & ~n742;
  assign n744 = ~n741 & ~n743;
  assign n745 = ~n742 & ~n743;
  assign n746 = ~n744 & ~n745;
  assign n747 = ~n633 & ~n638;
  assign n748 = ~n746 & ~n747;
  assign n749 = ~n746 & ~n748;
  assign n750 = ~n747 & ~n748;
  assign n751 = ~n749 & ~n750;
  assign n752 = 52 & 426;
  assign n753 = ~n751 & ~n752;
  assign n754 = ~n751 & ~n753;
  assign n755 = ~n752 & ~n753;
  assign n756 = ~n754 & ~n755;
  assign n757 = ~n643 & ~n648;
  assign n758 = ~n756 & ~n757;
  assign n759 = ~n756 & ~n758;
  assign n760 = ~n757 & ~n758;
  assign n761 = ~n759 & ~n760;
  assign n762 = 35 & 443;
  assign n763 = ~n761 & ~n762;
  assign n764 = ~n761 & ~n763;
  assign n765 = ~n762 & ~n763;
  assign n766 = ~n764 & ~n765;
  assign n767 = ~n653 & ~n658;
  assign n768 = ~n766 & ~n767;
  assign n769 = ~n766 & ~n768;
  assign n770 = ~n767 & ~n768;
  assign n771 = ~n769 & ~n770;
  assign n772 = 18 & 460;
  assign n773 = ~n771 & ~n772;
  assign n774 = ~n771 & ~n773;
  assign n775 = ~n772 & ~n773;
  assign n776 = ~n774 & ~n775;
  assign n777 = ~n663 & ~n668;
  assign n778 = ~n776 & ~n777;
  assign n779 = ~n776 & ~n778;
  assign n780 = ~n777 & ~n778;
  assign n781 = ~n779 & ~n780;
  assign n782 = \1  & 477;
  assign n783 = ~n781 & ~n782;
  assign n784 = ~n781 & ~n783;
  assign n785 = ~n782 & ~n783;
  assign 5308 = ~n784 & ~n785;
  assign n787 = 222 & 273;
  assign n788 = 205 & 290;
  assign n789 = n787 & ~n788;
  assign n790 = n787 & ~n789;
  assign n791 = ~n788 & ~n789;
  assign n792 = ~n790 & ~n791;
  assign n793 = ~n675 & ~n792;
  assign n794 = ~n792 & ~n793;
  assign n795 = ~n675 & ~n793;
  assign n796 = ~n794 & ~n795;
  assign n797 = 188 & 307;
  assign n798 = ~n796 & ~n797;
  assign n799 = ~n796 & ~n798;
  assign n800 = ~n797 & ~n798;
  assign n801 = ~n799 & ~n800;
  assign n802 = ~n678 & ~n683;
  assign n803 = ~n801 & ~n802;
  assign n804 = ~n801 & ~n803;
  assign n805 = ~n802 & ~n803;
  assign n806 = ~n804 & ~n805;
  assign n807 = 171 & 324;
  assign n808 = ~n806 & ~n807;
  assign n809 = ~n806 & ~n808;
  assign n810 = ~n807 & ~n808;
  assign n811 = ~n809 & ~n810;
  assign n812 = ~n688 & ~n693;
  assign n813 = ~n811 & ~n812;
  assign n814 = ~n811 & ~n813;
  assign n815 = ~n812 & ~n813;
  assign n816 = ~n814 & ~n815;
  assign n817 = 154 & 341;
  assign n818 = ~n816 & ~n817;
  assign n819 = ~n816 & ~n818;
  assign n820 = ~n817 & ~n818;
  assign n821 = ~n819 & ~n820;
  assign n822 = ~n698 & ~n703;
  assign n823 = ~n821 & ~n822;
  assign n824 = ~n821 & ~n823;
  assign n825 = ~n822 & ~n823;
  assign n826 = ~n824 & ~n825;
  assign n827 = 137 & 358;
  assign n828 = ~n826 & ~n827;
  assign n829 = ~n826 & ~n828;
  assign n830 = ~n827 & ~n828;
  assign n831 = ~n829 & ~n830;
  assign n832 = ~n708 & ~n713;
  assign n833 = ~n831 & ~n832;
  assign n834 = ~n831 & ~n833;
  assign n835 = ~n832 & ~n833;
  assign n836 = ~n834 & ~n835;
  assign n837 = 120 & 375;
  assign n838 = ~n836 & ~n837;
  assign n839 = ~n836 & ~n838;
  assign n840 = ~n837 & ~n838;
  assign n841 = ~n839 & ~n840;
  assign n842 = ~n718 & ~n723;
  assign n843 = ~n841 & ~n842;
  assign n844 = ~n841 & ~n843;
  assign n845 = ~n842 & ~n843;
  assign n846 = ~n844 & ~n845;
  assign n847 = 103 & 392;
  assign n848 = ~n846 & ~n847;
  assign n849 = ~n846 & ~n848;
  assign n850 = ~n847 & ~n848;
  assign n851 = ~n849 & ~n850;
  assign n852 = ~n728 & ~n733;
  assign n853 = ~n851 & ~n852;
  assign n854 = ~n851 & ~n853;
  assign n855 = ~n852 & ~n853;
  assign n856 = ~n854 & ~n855;
  assign n857 = 86 & 409;
  assign n858 = ~n856 & ~n857;
  assign n859 = ~n856 & ~n858;
  assign n860 = ~n857 & ~n858;
  assign n861 = ~n859 & ~n860;
  assign n862 = ~n738 & ~n743;
  assign n863 = ~n861 & ~n862;
  assign n864 = ~n861 & ~n863;
  assign n865 = ~n862 & ~n863;
  assign n866 = ~n864 & ~n865;
  assign n867 = 69 & 426;
  assign n868 = ~n866 & ~n867;
  assign n869 = ~n866 & ~n868;
  assign n870 = ~n867 & ~n868;
  assign n871 = ~n869 & ~n870;
  assign n872 = ~n748 & ~n753;
  assign n873 = ~n871 & ~n872;
  assign n874 = ~n871 & ~n873;
  assign n875 = ~n872 & ~n873;
  assign n876 = ~n874 & ~n875;
  assign n877 = 52 & 443;
  assign n878 = ~n876 & ~n877;
  assign n879 = ~n876 & ~n878;
  assign n880 = ~n877 & ~n878;
  assign n881 = ~n879 & ~n880;
  assign n882 = ~n758 & ~n763;
  assign n883 = ~n881 & ~n882;
  assign n884 = ~n881 & ~n883;
  assign n885 = ~n882 & ~n883;
  assign n886 = ~n884 & ~n885;
  assign n887 = 35 & 460;
  assign n888 = ~n886 & ~n887;
  assign n889 = ~n886 & ~n888;
  assign n890 = ~n887 & ~n888;
  assign n891 = ~n889 & ~n890;
  assign n892 = ~n768 & ~n773;
  assign n893 = ~n891 & ~n892;
  assign n894 = ~n891 & ~n893;
  assign n895 = ~n892 & ~n893;
  assign n896 = ~n894 & ~n895;
  assign n897 = 18 & 477;
  assign n898 = ~n896 & ~n897;
  assign n899 = ~n896 & ~n898;
  assign n900 = ~n897 & ~n898;
  assign n901 = ~n899 & ~n900;
  assign n902 = ~n778 & ~n783;
  assign n903 = ~n901 & ~n902;
  assign n904 = ~n901 & ~n903;
  assign n905 = ~n902 & ~n903;
  assign n906 = ~n904 & ~n905;
  assign n907 = \1  & 494;
  assign n908 = ~n906 & ~n907;
  assign n909 = ~n906 & ~n908;
  assign n910 = ~n907 & ~n908;
  assign 5672 = ~n909 & ~n910;
  assign n912 = 239 & 273;
  assign n913 = 222 & 290;
  assign n914 = n912 & ~n913;
  assign n915 = n912 & ~n914;
  assign n916 = ~n913 & ~n914;
  assign n917 = ~n915 & ~n916;
  assign n918 = ~n790 & ~n917;
  assign n919 = ~n917 & ~n918;
  assign n920 = ~n790 & ~n918;
  assign n921 = ~n919 & ~n920;
  assign n922 = 205 & 307;
  assign n923 = ~n921 & ~n922;
  assign n924 = ~n921 & ~n923;
  assign n925 = ~n922 & ~n923;
  assign n926 = ~n924 & ~n925;
  assign n927 = ~n793 & ~n798;
  assign n928 = ~n926 & ~n927;
  assign n929 = ~n926 & ~n928;
  assign n930 = ~n927 & ~n928;
  assign n931 = ~n929 & ~n930;
  assign n932 = 188 & 324;
  assign n933 = ~n931 & ~n932;
  assign n934 = ~n931 & ~n933;
  assign n935 = ~n932 & ~n933;
  assign n936 = ~n934 & ~n935;
  assign n937 = ~n803 & ~n808;
  assign n938 = ~n936 & ~n937;
  assign n939 = ~n936 & ~n938;
  assign n940 = ~n937 & ~n938;
  assign n941 = ~n939 & ~n940;
  assign n942 = 171 & 341;
  assign n943 = ~n941 & ~n942;
  assign n944 = ~n941 & ~n943;
  assign n945 = ~n942 & ~n943;
  assign n946 = ~n944 & ~n945;
  assign n947 = ~n813 & ~n818;
  assign n948 = ~n946 & ~n947;
  assign n949 = ~n946 & ~n948;
  assign n950 = ~n947 & ~n948;
  assign n951 = ~n949 & ~n950;
  assign n952 = 154 & 358;
  assign n953 = ~n951 & ~n952;
  assign n954 = ~n951 & ~n953;
  assign n955 = ~n952 & ~n953;
  assign n956 = ~n954 & ~n955;
  assign n957 = ~n823 & ~n828;
  assign n958 = ~n956 & ~n957;
  assign n959 = ~n956 & ~n958;
  assign n960 = ~n957 & ~n958;
  assign n961 = ~n959 & ~n960;
  assign n962 = 137 & 375;
  assign n963 = ~n961 & ~n962;
  assign n964 = ~n961 & ~n963;
  assign n965 = ~n962 & ~n963;
  assign n966 = ~n964 & ~n965;
  assign n967 = ~n833 & ~n838;
  assign n968 = ~n966 & ~n967;
  assign n969 = ~n966 & ~n968;
  assign n970 = ~n967 & ~n968;
  assign n971 = ~n969 & ~n970;
  assign n972 = 120 & 392;
  assign n973 = ~n971 & ~n972;
  assign n974 = ~n971 & ~n973;
  assign n975 = ~n972 & ~n973;
  assign n976 = ~n974 & ~n975;
  assign n977 = ~n843 & ~n848;
  assign n978 = ~n976 & ~n977;
  assign n979 = ~n976 & ~n978;
  assign n980 = ~n977 & ~n978;
  assign n981 = ~n979 & ~n980;
  assign n982 = 103 & 409;
  assign n983 = ~n981 & ~n982;
  assign n984 = ~n981 & ~n983;
  assign n985 = ~n982 & ~n983;
  assign n986 = ~n984 & ~n985;
  assign n987 = ~n853 & ~n858;
  assign n988 = ~n986 & ~n987;
  assign n989 = ~n986 & ~n988;
  assign n990 = ~n987 & ~n988;
  assign n991 = ~n989 & ~n990;
  assign n992 = 86 & 426;
  assign n993 = ~n991 & ~n992;
  assign n994 = ~n991 & ~n993;
  assign n995 = ~n992 & ~n993;
  assign n996 = ~n994 & ~n995;
  assign n997 = ~n863 & ~n868;
  assign n998 = ~n996 & ~n997;
  assign n999 = ~n996 & ~n998;
  assign n1000 = ~n997 & ~n998;
  assign n1001 = ~n999 & ~n1000;
  assign n1002 = 69 & 443;
  assign n1003 = ~n1001 & ~n1002;
  assign n1004 = ~n1001 & ~n1003;
  assign n1005 = ~n1002 & ~n1003;
  assign n1006 = ~n1004 & ~n1005;
  assign n1007 = ~n873 & ~n878;
  assign n1008 = ~n1006 & ~n1007;
  assign n1009 = ~n1006 & ~n1008;
  assign n1010 = ~n1007 & ~n1008;
  assign n1011 = ~n1009 & ~n1010;
  assign n1012 = 52 & 460;
  assign n1013 = ~n1011 & ~n1012;
  assign n1014 = ~n1011 & ~n1013;
  assign n1015 = ~n1012 & ~n1013;
  assign n1016 = ~n1014 & ~n1015;
  assign n1017 = ~n883 & ~n888;
  assign n1018 = ~n1016 & ~n1017;
  assign n1019 = ~n1016 & ~n1018;
  assign n1020 = ~n1017 & ~n1018;
  assign n1021 = ~n1019 & ~n1020;
  assign n1022 = 35 & 477;
  assign n1023 = ~n1021 & ~n1022;
  assign n1024 = ~n1021 & ~n1023;
  assign n1025 = ~n1022 & ~n1023;
  assign n1026 = ~n1024 & ~n1025;
  assign n1027 = ~n893 & ~n898;
  assign n1028 = ~n1026 & ~n1027;
  assign n1029 = ~n1026 & ~n1028;
  assign n1030 = ~n1027 & ~n1028;
  assign n1031 = ~n1029 & ~n1030;
  assign n1032 = 18 & 494;
  assign n1033 = ~n1031 & ~n1032;
  assign n1034 = ~n1031 & ~n1033;
  assign n1035 = ~n1032 & ~n1033;
  assign n1036 = ~n1034 & ~n1035;
  assign n1037 = ~n903 & ~n908;
  assign n1038 = ~n1036 & ~n1037;
  assign n1039 = ~n1036 & ~n1038;
  assign n1040 = ~n1037 & ~n1038;
  assign n1041 = ~n1039 & ~n1040;
  assign n1042 = \1  & 511;
  assign n1043 = ~n1041 & ~n1042;
  assign n1044 = ~n1041 & ~n1043;
  assign n1045 = ~n1042 & ~n1043;
  assign 5971 = ~n1044 & ~n1045;
  assign n1047 = 256 & 273;
  assign n1048 = 239 & 290;
  assign n1049 = n1047 & ~n1048;
  assign n1050 = n1047 & ~n1049;
  assign n1051 = ~n1048 & ~n1049;
  assign n1052 = ~n1050 & ~n1051;
  assign n1053 = ~n915 & ~n1052;
  assign n1054 = ~n1052 & ~n1053;
  assign n1055 = ~n915 & ~n1053;
  assign n1056 = ~n1054 & ~n1055;
  assign n1057 = 222 & 307;
  assign n1058 = ~n1056 & ~n1057;
  assign n1059 = ~n1056 & ~n1058;
  assign n1060 = ~n1057 & ~n1058;
  assign n1061 = ~n1059 & ~n1060;
  assign n1062 = ~n918 & ~n923;
  assign n1063 = ~n1061 & ~n1062;
  assign n1064 = ~n1061 & ~n1063;
  assign n1065 = ~n1062 & ~n1063;
  assign n1066 = ~n1064 & ~n1065;
  assign n1067 = 205 & 324;
  assign n1068 = ~n1066 & ~n1067;
  assign n1069 = ~n1066 & ~n1068;
  assign n1070 = ~n1067 & ~n1068;
  assign n1071 = ~n1069 & ~n1070;
  assign n1072 = ~n928 & ~n933;
  assign n1073 = ~n1071 & ~n1072;
  assign n1074 = ~n1071 & ~n1073;
  assign n1075 = ~n1072 & ~n1073;
  assign n1076 = ~n1074 & ~n1075;
  assign n1077 = 188 & 341;
  assign n1078 = ~n1076 & ~n1077;
  assign n1079 = ~n1076 & ~n1078;
  assign n1080 = ~n1077 & ~n1078;
  assign n1081 = ~n1079 & ~n1080;
  assign n1082 = ~n938 & ~n943;
  assign n1083 = ~n1081 & ~n1082;
  assign n1084 = ~n1081 & ~n1083;
  assign n1085 = ~n1082 & ~n1083;
  assign n1086 = ~n1084 & ~n1085;
  assign n1087 = 171 & 358;
  assign n1088 = ~n1086 & ~n1087;
  assign n1089 = ~n1086 & ~n1088;
  assign n1090 = ~n1087 & ~n1088;
  assign n1091 = ~n1089 & ~n1090;
  assign n1092 = ~n948 & ~n953;
  assign n1093 = ~n1091 & ~n1092;
  assign n1094 = ~n1091 & ~n1093;
  assign n1095 = ~n1092 & ~n1093;
  assign n1096 = ~n1094 & ~n1095;
  assign n1097 = 154 & 375;
  assign n1098 = ~n1096 & ~n1097;
  assign n1099 = ~n1096 & ~n1098;
  assign n1100 = ~n1097 & ~n1098;
  assign n1101 = ~n1099 & ~n1100;
  assign n1102 = ~n958 & ~n963;
  assign n1103 = ~n1101 & ~n1102;
  assign n1104 = ~n1101 & ~n1103;
  assign n1105 = ~n1102 & ~n1103;
  assign n1106 = ~n1104 & ~n1105;
  assign n1107 = 137 & 392;
  assign n1108 = ~n1106 & ~n1107;
  assign n1109 = ~n1106 & ~n1108;
  assign n1110 = ~n1107 & ~n1108;
  assign n1111 = ~n1109 & ~n1110;
  assign n1112 = ~n968 & ~n973;
  assign n1113 = ~n1111 & ~n1112;
  assign n1114 = ~n1111 & ~n1113;
  assign n1115 = ~n1112 & ~n1113;
  assign n1116 = ~n1114 & ~n1115;
  assign n1117 = 120 & 409;
  assign n1118 = ~n1116 & ~n1117;
  assign n1119 = ~n1116 & ~n1118;
  assign n1120 = ~n1117 & ~n1118;
  assign n1121 = ~n1119 & ~n1120;
  assign n1122 = ~n978 & ~n983;
  assign n1123 = ~n1121 & ~n1122;
  assign n1124 = ~n1121 & ~n1123;
  assign n1125 = ~n1122 & ~n1123;
  assign n1126 = ~n1124 & ~n1125;
  assign n1127 = 103 & 426;
  assign n1128 = ~n1126 & ~n1127;
  assign n1129 = ~n1126 & ~n1128;
  assign n1130 = ~n1127 & ~n1128;
  assign n1131 = ~n1129 & ~n1130;
  assign n1132 = ~n988 & ~n993;
  assign n1133 = ~n1131 & ~n1132;
  assign n1134 = ~n1131 & ~n1133;
  assign n1135 = ~n1132 & ~n1133;
  assign n1136 = ~n1134 & ~n1135;
  assign n1137 = 86 & 443;
  assign n1138 = ~n1136 & ~n1137;
  assign n1139 = ~n1136 & ~n1138;
  assign n1140 = ~n1137 & ~n1138;
  assign n1141 = ~n1139 & ~n1140;
  assign n1142 = ~n998 & ~n1003;
  assign n1143 = ~n1141 & ~n1142;
  assign n1144 = ~n1141 & ~n1143;
  assign n1145 = ~n1142 & ~n1143;
  assign n1146 = ~n1144 & ~n1145;
  assign n1147 = 69 & 460;
  assign n1148 = ~n1146 & ~n1147;
  assign n1149 = ~n1146 & ~n1148;
  assign n1150 = ~n1147 & ~n1148;
  assign n1151 = ~n1149 & ~n1150;
  assign n1152 = ~n1008 & ~n1013;
  assign n1153 = ~n1151 & ~n1152;
  assign n1154 = ~n1151 & ~n1153;
  assign n1155 = ~n1152 & ~n1153;
  assign n1156 = ~n1154 & ~n1155;
  assign n1157 = 52 & 477;
  assign n1158 = ~n1156 & ~n1157;
  assign n1159 = ~n1156 & ~n1158;
  assign n1160 = ~n1157 & ~n1158;
  assign n1161 = ~n1159 & ~n1160;
  assign n1162 = ~n1018 & ~n1023;
  assign n1163 = ~n1161 & ~n1162;
  assign n1164 = ~n1161 & ~n1163;
  assign n1165 = ~n1162 & ~n1163;
  assign n1166 = ~n1164 & ~n1165;
  assign n1167 = 35 & 494;
  assign n1168 = ~n1166 & ~n1167;
  assign n1169 = ~n1166 & ~n1168;
  assign n1170 = ~n1167 & ~n1168;
  assign n1171 = ~n1169 & ~n1170;
  assign n1172 = ~n1028 & ~n1033;
  assign n1173 = ~n1171 & ~n1172;
  assign n1174 = ~n1171 & ~n1173;
  assign n1175 = ~n1172 & ~n1173;
  assign n1176 = ~n1174 & ~n1175;
  assign n1177 = 18 & 511;
  assign n1178 = ~n1176 & ~n1177;
  assign n1179 = ~n1176 & ~n1178;
  assign n1180 = ~n1177 & ~n1178;
  assign n1181 = ~n1179 & ~n1180;
  assign n1182 = ~n1038 & ~n1043;
  assign n1183 = ~n1181 & ~n1182;
  assign n1184 = ~n1181 & ~n1183;
  assign n1185 = ~n1182 & ~n1183;
  assign n1186 = ~n1184 & ~n1185;
  assign n1187 = \1  & 528;
  assign n1188 = ~n1186 & ~n1187;
  assign n1189 = ~n1186 & ~n1188;
  assign n1190 = ~n1187 & ~n1188;
  assign 6123 = ~n1189 & ~n1190;
  assign n1192 = 256 & 290;
  assign n1193 = ~n1050 & ~n1192;
  assign n1194 = ~n1192 & ~n1193;
  assign n1195 = ~n1050 & ~n1193;
  assign n1196 = ~n1194 & ~n1195;
  assign n1197 = 239 & 307;
  assign n1198 = ~n1196 & ~n1197;
  assign n1199 = ~n1196 & ~n1198;
  assign n1200 = ~n1197 & ~n1198;
  assign n1201 = ~n1199 & ~n1200;
  assign n1202 = ~n1053 & ~n1058;
  assign n1203 = ~n1201 & ~n1202;
  assign n1204 = ~n1201 & ~n1203;
  assign n1205 = ~n1202 & ~n1203;
  assign n1206 = ~n1204 & ~n1205;
  assign n1207 = 222 & 324;
  assign n1208 = ~n1206 & ~n1207;
  assign n1209 = ~n1206 & ~n1208;
  assign n1210 = ~n1207 & ~n1208;
  assign n1211 = ~n1209 & ~n1210;
  assign n1212 = ~n1063 & ~n1068;
  assign n1213 = ~n1211 & ~n1212;
  assign n1214 = ~n1211 & ~n1213;
  assign n1215 = ~n1212 & ~n1213;
  assign n1216 = ~n1214 & ~n1215;
  assign n1217 = 205 & 341;
  assign n1218 = ~n1216 & ~n1217;
  assign n1219 = ~n1216 & ~n1218;
  assign n1220 = ~n1217 & ~n1218;
  assign n1221 = ~n1219 & ~n1220;
  assign n1222 = ~n1073 & ~n1078;
  assign n1223 = ~n1221 & ~n1222;
  assign n1224 = ~n1221 & ~n1223;
  assign n1225 = ~n1222 & ~n1223;
  assign n1226 = ~n1224 & ~n1225;
  assign n1227 = 188 & 358;
  assign n1228 = ~n1226 & ~n1227;
  assign n1229 = ~n1226 & ~n1228;
  assign n1230 = ~n1227 & ~n1228;
  assign n1231 = ~n1229 & ~n1230;
  assign n1232 = ~n1083 & ~n1088;
  assign n1233 = ~n1231 & ~n1232;
  assign n1234 = ~n1231 & ~n1233;
  assign n1235 = ~n1232 & ~n1233;
  assign n1236 = ~n1234 & ~n1235;
  assign n1237 = 171 & 375;
  assign n1238 = ~n1236 & ~n1237;
  assign n1239 = ~n1236 & ~n1238;
  assign n1240 = ~n1237 & ~n1238;
  assign n1241 = ~n1239 & ~n1240;
  assign n1242 = ~n1093 & ~n1098;
  assign n1243 = ~n1241 & ~n1242;
  assign n1244 = ~n1241 & ~n1243;
  assign n1245 = ~n1242 & ~n1243;
  assign n1246 = ~n1244 & ~n1245;
  assign n1247 = 154 & 392;
  assign n1248 = ~n1246 & ~n1247;
  assign n1249 = ~n1246 & ~n1248;
  assign n1250 = ~n1247 & ~n1248;
  assign n1251 = ~n1249 & ~n1250;
  assign n1252 = ~n1103 & ~n1108;
  assign n1253 = ~n1251 & ~n1252;
  assign n1254 = ~n1251 & ~n1253;
  assign n1255 = ~n1252 & ~n1253;
  assign n1256 = ~n1254 & ~n1255;
  assign n1257 = 137 & 409;
  assign n1258 = ~n1256 & ~n1257;
  assign n1259 = ~n1256 & ~n1258;
  assign n1260 = ~n1257 & ~n1258;
  assign n1261 = ~n1259 & ~n1260;
  assign n1262 = ~n1113 & ~n1118;
  assign n1263 = ~n1261 & ~n1262;
  assign n1264 = ~n1261 & ~n1263;
  assign n1265 = ~n1262 & ~n1263;
  assign n1266 = ~n1264 & ~n1265;
  assign n1267 = 120 & 426;
  assign n1268 = ~n1266 & ~n1267;
  assign n1269 = ~n1266 & ~n1268;
  assign n1270 = ~n1267 & ~n1268;
  assign n1271 = ~n1269 & ~n1270;
  assign n1272 = ~n1123 & ~n1128;
  assign n1273 = ~n1271 & ~n1272;
  assign n1274 = ~n1271 & ~n1273;
  assign n1275 = ~n1272 & ~n1273;
  assign n1276 = ~n1274 & ~n1275;
  assign n1277 = 103 & 443;
  assign n1278 = ~n1276 & ~n1277;
  assign n1279 = ~n1276 & ~n1278;
  assign n1280 = ~n1277 & ~n1278;
  assign n1281 = ~n1279 & ~n1280;
  assign n1282 = ~n1133 & ~n1138;
  assign n1283 = ~n1281 & ~n1282;
  assign n1284 = ~n1281 & ~n1283;
  assign n1285 = ~n1282 & ~n1283;
  assign n1286 = ~n1284 & ~n1285;
  assign n1287 = 86 & 460;
  assign n1288 = ~n1286 & ~n1287;
  assign n1289 = ~n1286 & ~n1288;
  assign n1290 = ~n1287 & ~n1288;
  assign n1291 = ~n1289 & ~n1290;
  assign n1292 = ~n1143 & ~n1148;
  assign n1293 = ~n1291 & ~n1292;
  assign n1294 = ~n1291 & ~n1293;
  assign n1295 = ~n1292 & ~n1293;
  assign n1296 = ~n1294 & ~n1295;
  assign n1297 = 69 & 477;
  assign n1298 = ~n1296 & ~n1297;
  assign n1299 = ~n1296 & ~n1298;
  assign n1300 = ~n1297 & ~n1298;
  assign n1301 = ~n1299 & ~n1300;
  assign n1302 = ~n1153 & ~n1158;
  assign n1303 = ~n1301 & ~n1302;
  assign n1304 = ~n1301 & ~n1303;
  assign n1305 = ~n1302 & ~n1303;
  assign n1306 = ~n1304 & ~n1305;
  assign n1307 = 52 & 494;
  assign n1308 = ~n1306 & ~n1307;
  assign n1309 = ~n1306 & ~n1308;
  assign n1310 = ~n1307 & ~n1308;
  assign n1311 = ~n1309 & ~n1310;
  assign n1312 = ~n1163 & ~n1168;
  assign n1313 = ~n1311 & ~n1312;
  assign n1314 = ~n1311 & ~n1313;
  assign n1315 = ~n1312 & ~n1313;
  assign n1316 = ~n1314 & ~n1315;
  assign n1317 = 35 & 511;
  assign n1318 = ~n1316 & ~n1317;
  assign n1319 = ~n1316 & ~n1318;
  assign n1320 = ~n1317 & ~n1318;
  assign n1321 = ~n1319 & ~n1320;
  assign n1322 = ~n1173 & ~n1178;
  assign n1323 = ~n1321 & ~n1322;
  assign n1324 = ~n1321 & ~n1323;
  assign n1325 = ~n1322 & ~n1323;
  assign n1326 = ~n1324 & ~n1325;
  assign n1327 = 18 & 528;
  assign n1328 = ~n1326 & ~n1327;
  assign n1329 = ~n1326 & ~n1328;
  assign n1330 = ~n1327 & ~n1328;
  assign n1331 = ~n1329 & ~n1330;
  assign n1332 = ~n1183 & ~n1188;
  assign n1333 = ~n1331 & ~n1332;
  assign n1334 = ~n1331 & ~n1333;
  assign n1335 = ~n1332 & ~n1333;
  assign 6150 = n1334 | n1335;
  assign n1337 = 256 & 307;
  assign n1338 = ~n1193 & ~n1198;
  assign n1339 = ~n1337 & ~n1338;
  assign n1340 = ~n1337 & ~n1339;
  assign n1341 = ~n1338 & ~n1339;
  assign n1342 = ~n1340 & ~n1341;
  assign n1343 = 239 & 324;
  assign n1344 = ~n1342 & ~n1343;
  assign n1345 = ~n1342 & ~n1344;
  assign n1346 = ~n1343 & ~n1344;
  assign n1347 = ~n1345 & ~n1346;
  assign n1348 = ~n1203 & ~n1208;
  assign n1349 = ~n1347 & ~n1348;
  assign n1350 = ~n1347 & ~n1349;
  assign n1351 = ~n1348 & ~n1349;
  assign n1352 = ~n1350 & ~n1351;
  assign n1353 = 222 & 341;
  assign n1354 = ~n1352 & ~n1353;
  assign n1355 = ~n1352 & ~n1354;
  assign n1356 = ~n1353 & ~n1354;
  assign n1357 = ~n1355 & ~n1356;
  assign n1358 = ~n1213 & ~n1218;
  assign n1359 = ~n1357 & ~n1358;
  assign n1360 = ~n1357 & ~n1359;
  assign n1361 = ~n1358 & ~n1359;
  assign n1362 = ~n1360 & ~n1361;
  assign n1363 = 205 & 358;
  assign n1364 = ~n1362 & ~n1363;
  assign n1365 = ~n1362 & ~n1364;
  assign n1366 = ~n1363 & ~n1364;
  assign n1367 = ~n1365 & ~n1366;
  assign n1368 = ~n1223 & ~n1228;
  assign n1369 = ~n1367 & ~n1368;
  assign n1370 = ~n1367 & ~n1369;
  assign n1371 = ~n1368 & ~n1369;
  assign n1372 = ~n1370 & ~n1371;
  assign n1373 = 188 & 375;
  assign n1374 = ~n1372 & ~n1373;
  assign n1375 = ~n1372 & ~n1374;
  assign n1376 = ~n1373 & ~n1374;
  assign n1377 = ~n1375 & ~n1376;
  assign n1378 = ~n1233 & ~n1238;
  assign n1379 = ~n1377 & ~n1378;
  assign n1380 = ~n1377 & ~n1379;
  assign n1381 = ~n1378 & ~n1379;
  assign n1382 = ~n1380 & ~n1381;
  assign n1383 = 171 & 392;
  assign n1384 = ~n1382 & ~n1383;
  assign n1385 = ~n1382 & ~n1384;
  assign n1386 = ~n1383 & ~n1384;
  assign n1387 = ~n1385 & ~n1386;
  assign n1388 = ~n1243 & ~n1248;
  assign n1389 = ~n1387 & ~n1388;
  assign n1390 = ~n1387 & ~n1389;
  assign n1391 = ~n1388 & ~n1389;
  assign n1392 = ~n1390 & ~n1391;
  assign n1393 = 154 & 409;
  assign n1394 = ~n1392 & ~n1393;
  assign n1395 = ~n1392 & ~n1394;
  assign n1396 = ~n1393 & ~n1394;
  assign n1397 = ~n1395 & ~n1396;
  assign n1398 = ~n1253 & ~n1258;
  assign n1399 = ~n1397 & ~n1398;
  assign n1400 = ~n1397 & ~n1399;
  assign n1401 = ~n1398 & ~n1399;
  assign n1402 = ~n1400 & ~n1401;
  assign n1403 = 137 & 426;
  assign n1404 = ~n1402 & ~n1403;
  assign n1405 = ~n1402 & ~n1404;
  assign n1406 = ~n1403 & ~n1404;
  assign n1407 = ~n1405 & ~n1406;
  assign n1408 = ~n1263 & ~n1268;
  assign n1409 = ~n1407 & ~n1408;
  assign n1410 = ~n1407 & ~n1409;
  assign n1411 = ~n1408 & ~n1409;
  assign n1412 = ~n1410 & ~n1411;
  assign n1413 = 120 & 443;
  assign n1414 = ~n1412 & ~n1413;
  assign n1415 = ~n1412 & ~n1414;
  assign n1416 = ~n1413 & ~n1414;
  assign n1417 = ~n1415 & ~n1416;
  assign n1418 = ~n1273 & ~n1278;
  assign n1419 = ~n1417 & ~n1418;
  assign n1420 = ~n1417 & ~n1419;
  assign n1421 = ~n1418 & ~n1419;
  assign n1422 = ~n1420 & ~n1421;
  assign n1423 = 103 & 460;
  assign n1424 = ~n1422 & ~n1423;
  assign n1425 = ~n1422 & ~n1424;
  assign n1426 = ~n1423 & ~n1424;
  assign n1427 = ~n1425 & ~n1426;
  assign n1428 = ~n1283 & ~n1288;
  assign n1429 = ~n1427 & ~n1428;
  assign n1430 = ~n1427 & ~n1429;
  assign n1431 = ~n1428 & ~n1429;
  assign n1432 = ~n1430 & ~n1431;
  assign n1433 = 86 & 477;
  assign n1434 = ~n1432 & ~n1433;
  assign n1435 = ~n1432 & ~n1434;
  assign n1436 = ~n1433 & ~n1434;
  assign n1437 = ~n1435 & ~n1436;
  assign n1438 = ~n1293 & ~n1298;
  assign n1439 = ~n1437 & ~n1438;
  assign n1440 = ~n1437 & ~n1439;
  assign n1441 = ~n1438 & ~n1439;
  assign n1442 = ~n1440 & ~n1441;
  assign n1443 = 69 & 494;
  assign n1444 = ~n1442 & ~n1443;
  assign n1445 = ~n1442 & ~n1444;
  assign n1446 = ~n1443 & ~n1444;
  assign n1447 = ~n1445 & ~n1446;
  assign n1448 = ~n1303 & ~n1308;
  assign n1449 = ~n1447 & ~n1448;
  assign n1450 = ~n1447 & ~n1449;
  assign n1451 = ~n1448 & ~n1449;
  assign n1452 = ~n1450 & ~n1451;
  assign n1453 = 52 & 511;
  assign n1454 = ~n1452 & ~n1453;
  assign n1455 = ~n1452 & ~n1454;
  assign n1456 = ~n1453 & ~n1454;
  assign n1457 = ~n1455 & ~n1456;
  assign n1458 = ~n1313 & ~n1318;
  assign n1459 = ~n1457 & ~n1458;
  assign n1460 = ~n1457 & ~n1459;
  assign n1461 = ~n1458 & ~n1459;
  assign n1462 = ~n1460 & ~n1461;
  assign n1463 = 35 & 528;
  assign n1464 = ~n1462 & ~n1463;
  assign n1465 = ~n1462 & ~n1464;
  assign n1466 = ~n1463 & ~n1464;
  assign n1467 = ~n1465 & ~n1466;
  assign n1468 = ~n1323 & ~n1328;
  assign n1469 = ~n1467 & ~n1468;
  assign n1470 = ~n1467 & ~n1469;
  assign n1471 = ~n1468 & ~n1469;
  assign n1472 = ~n1470 & ~n1471;
  assign n1473 = ~n1333 & ~6150;
  assign n1474 = ~n1472 & ~n1473;
  assign n1475 = ~n1472 & ~n1474;
  assign n1476 = ~n1473 & ~n1474;
  assign 6160 = ~n1475 & ~n1476;
  assign n1478 = 256 & 324;
  assign n1479 = ~n1339 & ~n1344;
  assign n1480 = ~n1478 & ~n1479;
  assign n1481 = ~n1478 & ~n1480;
  assign n1482 = ~n1479 & ~n1480;
  assign n1483 = ~n1481 & ~n1482;
  assign n1484 = 239 & 341;
  assign n1485 = ~n1483 & ~n1484;
  assign n1486 = ~n1483 & ~n1485;
  assign n1487 = ~n1484 & ~n1485;
  assign n1488 = ~n1486 & ~n1487;
  assign n1489 = ~n1349 & ~n1354;
  assign n1490 = ~n1488 & ~n1489;
  assign n1491 = ~n1488 & ~n1490;
  assign n1492 = ~n1489 & ~n1490;
  assign n1493 = ~n1491 & ~n1492;
  assign n1494 = 222 & 358;
  assign n1495 = ~n1493 & ~n1494;
  assign n1496 = ~n1493 & ~n1495;
  assign n1497 = ~n1494 & ~n1495;
  assign n1498 = ~n1496 & ~n1497;
  assign n1499 = ~n1359 & ~n1364;
  assign n1500 = ~n1498 & ~n1499;
  assign n1501 = ~n1498 & ~n1500;
  assign n1502 = ~n1499 & ~n1500;
  assign n1503 = ~n1501 & ~n1502;
  assign n1504 = 205 & 375;
  assign n1505 = ~n1503 & ~n1504;
  assign n1506 = ~n1503 & ~n1505;
  assign n1507 = ~n1504 & ~n1505;
  assign n1508 = ~n1506 & ~n1507;
  assign n1509 = ~n1369 & ~n1374;
  assign n1510 = ~n1508 & ~n1509;
  assign n1511 = ~n1508 & ~n1510;
  assign n1512 = ~n1509 & ~n1510;
  assign n1513 = ~n1511 & ~n1512;
  assign n1514 = 188 & 392;
  assign n1515 = ~n1513 & ~n1514;
  assign n1516 = ~n1513 & ~n1515;
  assign n1517 = ~n1514 & ~n1515;
  assign n1518 = ~n1516 & ~n1517;
  assign n1519 = ~n1379 & ~n1384;
  assign n1520 = ~n1518 & ~n1519;
  assign n1521 = ~n1518 & ~n1520;
  assign n1522 = ~n1519 & ~n1520;
  assign n1523 = ~n1521 & ~n1522;
  assign n1524 = 171 & 409;
  assign n1525 = ~n1523 & ~n1524;
  assign n1526 = ~n1523 & ~n1525;
  assign n1527 = ~n1524 & ~n1525;
  assign n1528 = ~n1526 & ~n1527;
  assign n1529 = ~n1389 & ~n1394;
  assign n1530 = ~n1528 & ~n1529;
  assign n1531 = ~n1528 & ~n1530;
  assign n1532 = ~n1529 & ~n1530;
  assign n1533 = ~n1531 & ~n1532;
  assign n1534 = 154 & 426;
  assign n1535 = ~n1533 & ~n1534;
  assign n1536 = ~n1533 & ~n1535;
  assign n1537 = ~n1534 & ~n1535;
  assign n1538 = ~n1536 & ~n1537;
  assign n1539 = ~n1399 & ~n1404;
  assign n1540 = ~n1538 & ~n1539;
  assign n1541 = ~n1538 & ~n1540;
  assign n1542 = ~n1539 & ~n1540;
  assign n1543 = ~n1541 & ~n1542;
  assign n1544 = 137 & 443;
  assign n1545 = ~n1543 & ~n1544;
  assign n1546 = ~n1543 & ~n1545;
  assign n1547 = ~n1544 & ~n1545;
  assign n1548 = ~n1546 & ~n1547;
  assign n1549 = ~n1409 & ~n1414;
  assign n1550 = ~n1548 & ~n1549;
  assign n1551 = ~n1548 & ~n1550;
  assign n1552 = ~n1549 & ~n1550;
  assign n1553 = ~n1551 & ~n1552;
  assign n1554 = 120 & 460;
  assign n1555 = ~n1553 & ~n1554;
  assign n1556 = ~n1553 & ~n1555;
  assign n1557 = ~n1554 & ~n1555;
  assign n1558 = ~n1556 & ~n1557;
  assign n1559 = ~n1419 & ~n1424;
  assign n1560 = ~n1558 & ~n1559;
  assign n1561 = ~n1558 & ~n1560;
  assign n1562 = ~n1559 & ~n1560;
  assign n1563 = ~n1561 & ~n1562;
  assign n1564 = 103 & 477;
  assign n1565 = ~n1563 & ~n1564;
  assign n1566 = ~n1563 & ~n1565;
  assign n1567 = ~n1564 & ~n1565;
  assign n1568 = ~n1566 & ~n1567;
  assign n1569 = ~n1429 & ~n1434;
  assign n1570 = ~n1568 & ~n1569;
  assign n1571 = ~n1568 & ~n1570;
  assign n1572 = ~n1569 & ~n1570;
  assign n1573 = ~n1571 & ~n1572;
  assign n1574 = 86 & 494;
  assign n1575 = ~n1573 & ~n1574;
  assign n1576 = ~n1573 & ~n1575;
  assign n1577 = ~n1574 & ~n1575;
  assign n1578 = ~n1576 & ~n1577;
  assign n1579 = ~n1439 & ~n1444;
  assign n1580 = ~n1578 & ~n1579;
  assign n1581 = ~n1578 & ~n1580;
  assign n1582 = ~n1579 & ~n1580;
  assign n1583 = ~n1581 & ~n1582;
  assign n1584 = 69 & 511;
  assign n1585 = ~n1583 & ~n1584;
  assign n1586 = ~n1583 & ~n1585;
  assign n1587 = ~n1584 & ~n1585;
  assign n1588 = ~n1586 & ~n1587;
  assign n1589 = ~n1449 & ~n1454;
  assign n1590 = ~n1588 & ~n1589;
  assign n1591 = ~n1588 & ~n1590;
  assign n1592 = ~n1589 & ~n1590;
  assign n1593 = ~n1591 & ~n1592;
  assign n1594 = 52 & 528;
  assign n1595 = ~n1593 & ~n1594;
  assign n1596 = ~n1593 & ~n1595;
  assign n1597 = ~n1594 & ~n1595;
  assign n1598 = ~n1596 & ~n1597;
  assign n1599 = ~n1459 & ~n1464;
  assign n1600 = ~n1598 & ~n1599;
  assign n1601 = ~n1598 & ~n1600;
  assign n1602 = ~n1599 & ~n1600;
  assign n1603 = ~n1601 & ~n1602;
  assign n1604 = ~n1469 & ~n1474;
  assign n1605 = ~n1603 & ~n1604;
  assign n1606 = ~n1603 & ~n1605;
  assign n1607 = ~n1604 & ~n1605;
  assign 6170 = ~n1606 & ~n1607;
  assign n1609 = 256 & 341;
  assign n1610 = ~n1480 & ~n1485;
  assign n1611 = ~n1609 & ~n1610;
  assign n1612 = ~n1609 & ~n1611;
  assign n1613 = ~n1610 & ~n1611;
  assign n1614 = ~n1612 & ~n1613;
  assign n1615 = 239 & 358;
  assign n1616 = ~n1614 & ~n1615;
  assign n1617 = ~n1614 & ~n1616;
  assign n1618 = ~n1615 & ~n1616;
  assign n1619 = ~n1617 & ~n1618;
  assign n1620 = ~n1490 & ~n1495;
  assign n1621 = ~n1619 & ~n1620;
  assign n1622 = ~n1619 & ~n1621;
  assign n1623 = ~n1620 & ~n1621;
  assign n1624 = ~n1622 & ~n1623;
  assign n1625 = 222 & 375;
  assign n1626 = ~n1624 & ~n1625;
  assign n1627 = ~n1624 & ~n1626;
  assign n1628 = ~n1625 & ~n1626;
  assign n1629 = ~n1627 & ~n1628;
  assign n1630 = ~n1500 & ~n1505;
  assign n1631 = ~n1629 & ~n1630;
  assign n1632 = ~n1629 & ~n1631;
  assign n1633 = ~n1630 & ~n1631;
  assign n1634 = ~n1632 & ~n1633;
  assign n1635 = 205 & 392;
  assign n1636 = ~n1634 & ~n1635;
  assign n1637 = ~n1634 & ~n1636;
  assign n1638 = ~n1635 & ~n1636;
  assign n1639 = ~n1637 & ~n1638;
  assign n1640 = ~n1510 & ~n1515;
  assign n1641 = ~n1639 & ~n1640;
  assign n1642 = ~n1639 & ~n1641;
  assign n1643 = ~n1640 & ~n1641;
  assign n1644 = ~n1642 & ~n1643;
  assign n1645 = 188 & 409;
  assign n1646 = ~n1644 & ~n1645;
  assign n1647 = ~n1644 & ~n1646;
  assign n1648 = ~n1645 & ~n1646;
  assign n1649 = ~n1647 & ~n1648;
  assign n1650 = ~n1520 & ~n1525;
  assign n1651 = ~n1649 & ~n1650;
  assign n1652 = ~n1649 & ~n1651;
  assign n1653 = ~n1650 & ~n1651;
  assign n1654 = ~n1652 & ~n1653;
  assign n1655 = 171 & 426;
  assign n1656 = ~n1654 & ~n1655;
  assign n1657 = ~n1654 & ~n1656;
  assign n1658 = ~n1655 & ~n1656;
  assign n1659 = ~n1657 & ~n1658;
  assign n1660 = ~n1530 & ~n1535;
  assign n1661 = ~n1659 & ~n1660;
  assign n1662 = ~n1659 & ~n1661;
  assign n1663 = ~n1660 & ~n1661;
  assign n1664 = ~n1662 & ~n1663;
  assign n1665 = 154 & 443;
  assign n1666 = ~n1664 & ~n1665;
  assign n1667 = ~n1664 & ~n1666;
  assign n1668 = ~n1665 & ~n1666;
  assign n1669 = ~n1667 & ~n1668;
  assign n1670 = ~n1540 & ~n1545;
  assign n1671 = ~n1669 & ~n1670;
  assign n1672 = ~n1669 & ~n1671;
  assign n1673 = ~n1670 & ~n1671;
  assign n1674 = ~n1672 & ~n1673;
  assign n1675 = 137 & 460;
  assign n1676 = ~n1674 & ~n1675;
  assign n1677 = ~n1674 & ~n1676;
  assign n1678 = ~n1675 & ~n1676;
  assign n1679 = ~n1677 & ~n1678;
  assign n1680 = ~n1550 & ~n1555;
  assign n1681 = ~n1679 & ~n1680;
  assign n1682 = ~n1679 & ~n1681;
  assign n1683 = ~n1680 & ~n1681;
  assign n1684 = ~n1682 & ~n1683;
  assign n1685 = 120 & 477;
  assign n1686 = ~n1684 & ~n1685;
  assign n1687 = ~n1684 & ~n1686;
  assign n1688 = ~n1685 & ~n1686;
  assign n1689 = ~n1687 & ~n1688;
  assign n1690 = ~n1560 & ~n1565;
  assign n1691 = ~n1689 & ~n1690;
  assign n1692 = ~n1689 & ~n1691;
  assign n1693 = ~n1690 & ~n1691;
  assign n1694 = ~n1692 & ~n1693;
  assign n1695 = 103 & 494;
  assign n1696 = ~n1694 & ~n1695;
  assign n1697 = ~n1694 & ~n1696;
  assign n1698 = ~n1695 & ~n1696;
  assign n1699 = ~n1697 & ~n1698;
  assign n1700 = ~n1570 & ~n1575;
  assign n1701 = ~n1699 & ~n1700;
  assign n1702 = ~n1699 & ~n1701;
  assign n1703 = ~n1700 & ~n1701;
  assign n1704 = ~n1702 & ~n1703;
  assign n1705 = 86 & 511;
  assign n1706 = ~n1704 & ~n1705;
  assign n1707 = ~n1704 & ~n1706;
  assign n1708 = ~n1705 & ~n1706;
  assign n1709 = ~n1707 & ~n1708;
  assign n1710 = ~n1580 & ~n1585;
  assign n1711 = ~n1709 & ~n1710;
  assign n1712 = ~n1709 & ~n1711;
  assign n1713 = ~n1710 & ~n1711;
  assign n1714 = ~n1712 & ~n1713;
  assign n1715 = 69 & 528;
  assign n1716 = ~n1714 & ~n1715;
  assign n1717 = ~n1714 & ~n1716;
  assign n1718 = ~n1715 & ~n1716;
  assign n1719 = ~n1717 & ~n1718;
  assign n1720 = ~n1590 & ~n1595;
  assign n1721 = ~n1719 & ~n1720;
  assign n1722 = ~n1719 & ~n1721;
  assign n1723 = ~n1720 & ~n1721;
  assign n1724 = ~n1722 & ~n1723;
  assign n1725 = ~n1600 & ~n1605;
  assign n1726 = ~n1724 & ~n1725;
  assign n1727 = ~n1724 & ~n1726;
  assign n1728 = ~n1725 & ~n1726;
  assign 6180 = ~n1727 & ~n1728;
  assign n1730 = 256 & 358;
  assign n1731 = ~n1611 & ~n1616;
  assign n1732 = ~n1730 & ~n1731;
  assign n1733 = ~n1730 & ~n1732;
  assign n1734 = ~n1731 & ~n1732;
  assign n1735 = ~n1733 & ~n1734;
  assign n1736 = 239 & 375;
  assign n1737 = ~n1735 & ~n1736;
  assign n1738 = ~n1735 & ~n1737;
  assign n1739 = ~n1736 & ~n1737;
  assign n1740 = ~n1738 & ~n1739;
  assign n1741 = ~n1621 & ~n1626;
  assign n1742 = ~n1740 & ~n1741;
  assign n1743 = ~n1740 & ~n1742;
  assign n1744 = ~n1741 & ~n1742;
  assign n1745 = ~n1743 & ~n1744;
  assign n1746 = 222 & 392;
  assign n1747 = ~n1745 & ~n1746;
  assign n1748 = ~n1745 & ~n1747;
  assign n1749 = ~n1746 & ~n1747;
  assign n1750 = ~n1748 & ~n1749;
  assign n1751 = ~n1631 & ~n1636;
  assign n1752 = ~n1750 & ~n1751;
  assign n1753 = ~n1750 & ~n1752;
  assign n1754 = ~n1751 & ~n1752;
  assign n1755 = ~n1753 & ~n1754;
  assign n1756 = 205 & 409;
  assign n1757 = ~n1755 & ~n1756;
  assign n1758 = ~n1755 & ~n1757;
  assign n1759 = ~n1756 & ~n1757;
  assign n1760 = ~n1758 & ~n1759;
  assign n1761 = ~n1641 & ~n1646;
  assign n1762 = ~n1760 & ~n1761;
  assign n1763 = ~n1760 & ~n1762;
  assign n1764 = ~n1761 & ~n1762;
  assign n1765 = ~n1763 & ~n1764;
  assign n1766 = 188 & 426;
  assign n1767 = ~n1765 & ~n1766;
  assign n1768 = ~n1765 & ~n1767;
  assign n1769 = ~n1766 & ~n1767;
  assign n1770 = ~n1768 & ~n1769;
  assign n1771 = ~n1651 & ~n1656;
  assign n1772 = ~n1770 & ~n1771;
  assign n1773 = ~n1770 & ~n1772;
  assign n1774 = ~n1771 & ~n1772;
  assign n1775 = ~n1773 & ~n1774;
  assign n1776 = 171 & 443;
  assign n1777 = ~n1775 & ~n1776;
  assign n1778 = ~n1775 & ~n1777;
  assign n1779 = ~n1776 & ~n1777;
  assign n1780 = ~n1778 & ~n1779;
  assign n1781 = ~n1661 & ~n1666;
  assign n1782 = ~n1780 & ~n1781;
  assign n1783 = ~n1780 & ~n1782;
  assign n1784 = ~n1781 & ~n1782;
  assign n1785 = ~n1783 & ~n1784;
  assign n1786 = 154 & 460;
  assign n1787 = ~n1785 & ~n1786;
  assign n1788 = ~n1785 & ~n1787;
  assign n1789 = ~n1786 & ~n1787;
  assign n1790 = ~n1788 & ~n1789;
  assign n1791 = ~n1671 & ~n1676;
  assign n1792 = ~n1790 & ~n1791;
  assign n1793 = ~n1790 & ~n1792;
  assign n1794 = ~n1791 & ~n1792;
  assign n1795 = ~n1793 & ~n1794;
  assign n1796 = 137 & 477;
  assign n1797 = ~n1795 & ~n1796;
  assign n1798 = ~n1795 & ~n1797;
  assign n1799 = ~n1796 & ~n1797;
  assign n1800 = ~n1798 & ~n1799;
  assign n1801 = ~n1681 & ~n1686;
  assign n1802 = ~n1800 & ~n1801;
  assign n1803 = ~n1800 & ~n1802;
  assign n1804 = ~n1801 & ~n1802;
  assign n1805 = ~n1803 & ~n1804;
  assign n1806 = 120 & 494;
  assign n1807 = ~n1805 & ~n1806;
  assign n1808 = ~n1805 & ~n1807;
  assign n1809 = ~n1806 & ~n1807;
  assign n1810 = ~n1808 & ~n1809;
  assign n1811 = ~n1691 & ~n1696;
  assign n1812 = ~n1810 & ~n1811;
  assign n1813 = ~n1810 & ~n1812;
  assign n1814 = ~n1811 & ~n1812;
  assign n1815 = ~n1813 & ~n1814;
  assign n1816 = 103 & 511;
  assign n1817 = ~n1815 & ~n1816;
  assign n1818 = ~n1815 & ~n1817;
  assign n1819 = ~n1816 & ~n1817;
  assign n1820 = ~n1818 & ~n1819;
  assign n1821 = ~n1701 & ~n1706;
  assign n1822 = ~n1820 & ~n1821;
  assign n1823 = ~n1820 & ~n1822;
  assign n1824 = ~n1821 & ~n1822;
  assign n1825 = ~n1823 & ~n1824;
  assign n1826 = 86 & 528;
  assign n1827 = ~n1825 & ~n1826;
  assign n1828 = ~n1825 & ~n1827;
  assign n1829 = ~n1826 & ~n1827;
  assign n1830 = ~n1828 & ~n1829;
  assign n1831 = ~n1711 & ~n1716;
  assign n1832 = ~n1830 & ~n1831;
  assign n1833 = ~n1830 & ~n1832;
  assign n1834 = ~n1831 & ~n1832;
  assign n1835 = ~n1833 & ~n1834;
  assign n1836 = ~n1721 & ~n1726;
  assign n1837 = ~n1835 & ~n1836;
  assign n1838 = ~n1835 & ~n1837;
  assign n1839 = ~n1836 & ~n1837;
  assign 6190 = ~n1838 & ~n1839;
  assign n1841 = 256 & 375;
  assign n1842 = ~n1732 & ~n1737;
  assign n1843 = ~n1841 & ~n1842;
  assign n1844 = ~n1841 & ~n1843;
  assign n1845 = ~n1842 & ~n1843;
  assign n1846 = ~n1844 & ~n1845;
  assign n1847 = 239 & 392;
  assign n1848 = ~n1846 & ~n1847;
  assign n1849 = ~n1846 & ~n1848;
  assign n1850 = ~n1847 & ~n1848;
  assign n1851 = ~n1849 & ~n1850;
  assign n1852 = ~n1742 & ~n1747;
  assign n1853 = ~n1851 & ~n1852;
  assign n1854 = ~n1851 & ~n1853;
  assign n1855 = ~n1852 & ~n1853;
  assign n1856 = ~n1854 & ~n1855;
  assign n1857 = 222 & 409;
  assign n1858 = ~n1856 & ~n1857;
  assign n1859 = ~n1856 & ~n1858;
  assign n1860 = ~n1857 & ~n1858;
  assign n1861 = ~n1859 & ~n1860;
  assign n1862 = ~n1752 & ~n1757;
  assign n1863 = ~n1861 & ~n1862;
  assign n1864 = ~n1861 & ~n1863;
  assign n1865 = ~n1862 & ~n1863;
  assign n1866 = ~n1864 & ~n1865;
  assign n1867 = 205 & 426;
  assign n1868 = ~n1866 & ~n1867;
  assign n1869 = ~n1866 & ~n1868;
  assign n1870 = ~n1867 & ~n1868;
  assign n1871 = ~n1869 & ~n1870;
  assign n1872 = ~n1762 & ~n1767;
  assign n1873 = ~n1871 & ~n1872;
  assign n1874 = ~n1871 & ~n1873;
  assign n1875 = ~n1872 & ~n1873;
  assign n1876 = ~n1874 & ~n1875;
  assign n1877 = 188 & 443;
  assign n1878 = ~n1876 & ~n1877;
  assign n1879 = ~n1876 & ~n1878;
  assign n1880 = ~n1877 & ~n1878;
  assign n1881 = ~n1879 & ~n1880;
  assign n1882 = ~n1772 & ~n1777;
  assign n1883 = ~n1881 & ~n1882;
  assign n1884 = ~n1881 & ~n1883;
  assign n1885 = ~n1882 & ~n1883;
  assign n1886 = ~n1884 & ~n1885;
  assign n1887 = 171 & 460;
  assign n1888 = ~n1886 & ~n1887;
  assign n1889 = ~n1886 & ~n1888;
  assign n1890 = ~n1887 & ~n1888;
  assign n1891 = ~n1889 & ~n1890;
  assign n1892 = ~n1782 & ~n1787;
  assign n1893 = ~n1891 & ~n1892;
  assign n1894 = ~n1891 & ~n1893;
  assign n1895 = ~n1892 & ~n1893;
  assign n1896 = ~n1894 & ~n1895;
  assign n1897 = 154 & 477;
  assign n1898 = ~n1896 & ~n1897;
  assign n1899 = ~n1896 & ~n1898;
  assign n1900 = ~n1897 & ~n1898;
  assign n1901 = ~n1899 & ~n1900;
  assign n1902 = ~n1792 & ~n1797;
  assign n1903 = ~n1901 & ~n1902;
  assign n1904 = ~n1901 & ~n1903;
  assign n1905 = ~n1902 & ~n1903;
  assign n1906 = ~n1904 & ~n1905;
  assign n1907 = 137 & 494;
  assign n1908 = ~n1906 & ~n1907;
  assign n1909 = ~n1906 & ~n1908;
  assign n1910 = ~n1907 & ~n1908;
  assign n1911 = ~n1909 & ~n1910;
  assign n1912 = ~n1802 & ~n1807;
  assign n1913 = ~n1911 & ~n1912;
  assign n1914 = ~n1911 & ~n1913;
  assign n1915 = ~n1912 & ~n1913;
  assign n1916 = ~n1914 & ~n1915;
  assign n1917 = 120 & 511;
  assign n1918 = ~n1916 & ~n1917;
  assign n1919 = ~n1916 & ~n1918;
  assign n1920 = ~n1917 & ~n1918;
  assign n1921 = ~n1919 & ~n1920;
  assign n1922 = ~n1812 & ~n1817;
  assign n1923 = ~n1921 & ~n1922;
  assign n1924 = ~n1921 & ~n1923;
  assign n1925 = ~n1922 & ~n1923;
  assign n1926 = ~n1924 & ~n1925;
  assign n1927 = 103 & 528;
  assign n1928 = ~n1926 & ~n1927;
  assign n1929 = ~n1926 & ~n1928;
  assign n1930 = ~n1927 & ~n1928;
  assign n1931 = ~n1929 & ~n1930;
  assign n1932 = ~n1822 & ~n1827;
  assign n1933 = ~n1931 & ~n1932;
  assign n1934 = ~n1931 & ~n1933;
  assign n1935 = ~n1932 & ~n1933;
  assign n1936 = ~n1934 & ~n1935;
  assign n1937 = ~n1832 & ~n1837;
  assign n1938 = ~n1936 & ~n1937;
  assign n1939 = ~n1936 & ~n1938;
  assign n1940 = ~n1937 & ~n1938;
  assign 6200 = ~n1939 & ~n1940;
  assign n1942 = 256 & 392;
  assign n1943 = ~n1843 & ~n1848;
  assign n1944 = ~n1942 & ~n1943;
  assign n1945 = ~n1942 & ~n1944;
  assign n1946 = ~n1943 & ~n1944;
  assign n1947 = ~n1945 & ~n1946;
  assign n1948 = 239 & 409;
  assign n1949 = ~n1947 & ~n1948;
  assign n1950 = ~n1947 & ~n1949;
  assign n1951 = ~n1948 & ~n1949;
  assign n1952 = ~n1950 & ~n1951;
  assign n1953 = ~n1853 & ~n1858;
  assign n1954 = ~n1952 & ~n1953;
  assign n1955 = ~n1952 & ~n1954;
  assign n1956 = ~n1953 & ~n1954;
  assign n1957 = ~n1955 & ~n1956;
  assign n1958 = 222 & 426;
  assign n1959 = ~n1957 & ~n1958;
  assign n1960 = ~n1957 & ~n1959;
  assign n1961 = ~n1958 & ~n1959;
  assign n1962 = ~n1960 & ~n1961;
  assign n1963 = ~n1863 & ~n1868;
  assign n1964 = ~n1962 & ~n1963;
  assign n1965 = ~n1962 & ~n1964;
  assign n1966 = ~n1963 & ~n1964;
  assign n1967 = ~n1965 & ~n1966;
  assign n1968 = 205 & 443;
  assign n1969 = ~n1967 & ~n1968;
  assign n1970 = ~n1967 & ~n1969;
  assign n1971 = ~n1968 & ~n1969;
  assign n1972 = ~n1970 & ~n1971;
  assign n1973 = ~n1873 & ~n1878;
  assign n1974 = ~n1972 & ~n1973;
  assign n1975 = ~n1972 & ~n1974;
  assign n1976 = ~n1973 & ~n1974;
  assign n1977 = ~n1975 & ~n1976;
  assign n1978 = 188 & 460;
  assign n1979 = ~n1977 & ~n1978;
  assign n1980 = ~n1977 & ~n1979;
  assign n1981 = ~n1978 & ~n1979;
  assign n1982 = ~n1980 & ~n1981;
  assign n1983 = ~n1883 & ~n1888;
  assign n1984 = ~n1982 & ~n1983;
  assign n1985 = ~n1982 & ~n1984;
  assign n1986 = ~n1983 & ~n1984;
  assign n1987 = ~n1985 & ~n1986;
  assign n1988 = 171 & 477;
  assign n1989 = ~n1987 & ~n1988;
  assign n1990 = ~n1987 & ~n1989;
  assign n1991 = ~n1988 & ~n1989;
  assign n1992 = ~n1990 & ~n1991;
  assign n1993 = ~n1893 & ~n1898;
  assign n1994 = ~n1992 & ~n1993;
  assign n1995 = ~n1992 & ~n1994;
  assign n1996 = ~n1993 & ~n1994;
  assign n1997 = ~n1995 & ~n1996;
  assign n1998 = 154 & 494;
  assign n1999 = ~n1997 & ~n1998;
  assign n2000 = ~n1997 & ~n1999;
  assign n2001 = ~n1998 & ~n1999;
  assign n2002 = ~n2000 & ~n2001;
  assign n2003 = ~n1903 & ~n1908;
  assign n2004 = ~n2002 & ~n2003;
  assign n2005 = ~n2002 & ~n2004;
  assign n2006 = ~n2003 & ~n2004;
  assign n2007 = ~n2005 & ~n2006;
  assign n2008 = 137 & 511;
  assign n2009 = ~n2007 & ~n2008;
  assign n2010 = ~n2007 & ~n2009;
  assign n2011 = ~n2008 & ~n2009;
  assign n2012 = ~n2010 & ~n2011;
  assign n2013 = ~n1913 & ~n1918;
  assign n2014 = ~n2012 & ~n2013;
  assign n2015 = ~n2012 & ~n2014;
  assign n2016 = ~n2013 & ~n2014;
  assign n2017 = ~n2015 & ~n2016;
  assign n2018 = 120 & 528;
  assign n2019 = ~n2017 & ~n2018;
  assign n2020 = ~n2017 & ~n2019;
  assign n2021 = ~n2018 & ~n2019;
  assign n2022 = ~n2020 & ~n2021;
  assign n2023 = ~n1923 & ~n1928;
  assign n2024 = ~n2022 & ~n2023;
  assign n2025 = ~n2022 & ~n2024;
  assign n2026 = ~n2023 & ~n2024;
  assign n2027 = ~n2025 & ~n2026;
  assign n2028 = ~n1933 & ~n1938;
  assign n2029 = ~n2027 & ~n2028;
  assign n2030 = ~n2027 & ~n2029;
  assign n2031 = ~n2028 & ~n2029;
  assign 6210 = ~n2030 & ~n2031;
  assign n2033 = 256 & 409;
  assign n2034 = ~n1944 & ~n1949;
  assign n2035 = ~n2033 & ~n2034;
  assign n2036 = ~n2033 & ~n2035;
  assign n2037 = ~n2034 & ~n2035;
  assign n2038 = ~n2036 & ~n2037;
  assign n2039 = 239 & 426;
  assign n2040 = ~n2038 & ~n2039;
  assign n2041 = ~n2038 & ~n2040;
  assign n2042 = ~n2039 & ~n2040;
  assign n2043 = ~n2041 & ~n2042;
  assign n2044 = ~n1954 & ~n1959;
  assign n2045 = ~n2043 & ~n2044;
  assign n2046 = ~n2043 & ~n2045;
  assign n2047 = ~n2044 & ~n2045;
  assign n2048 = ~n2046 & ~n2047;
  assign n2049 = 222 & 443;
  assign n2050 = ~n2048 & ~n2049;
  assign n2051 = ~n2048 & ~n2050;
  assign n2052 = ~n2049 & ~n2050;
  assign n2053 = ~n2051 & ~n2052;
  assign n2054 = ~n1964 & ~n1969;
  assign n2055 = ~n2053 & ~n2054;
  assign n2056 = ~n2053 & ~n2055;
  assign n2057 = ~n2054 & ~n2055;
  assign n2058 = ~n2056 & ~n2057;
  assign n2059 = 205 & 460;
  assign n2060 = ~n2058 & ~n2059;
  assign n2061 = ~n2058 & ~n2060;
  assign n2062 = ~n2059 & ~n2060;
  assign n2063 = ~n2061 & ~n2062;
  assign n2064 = ~n1974 & ~n1979;
  assign n2065 = ~n2063 & ~n2064;
  assign n2066 = ~n2063 & ~n2065;
  assign n2067 = ~n2064 & ~n2065;
  assign n2068 = ~n2066 & ~n2067;
  assign n2069 = 188 & 477;
  assign n2070 = ~n2068 & ~n2069;
  assign n2071 = ~n2068 & ~n2070;
  assign n2072 = ~n2069 & ~n2070;
  assign n2073 = ~n2071 & ~n2072;
  assign n2074 = ~n1984 & ~n1989;
  assign n2075 = ~n2073 & ~n2074;
  assign n2076 = ~n2073 & ~n2075;
  assign n2077 = ~n2074 & ~n2075;
  assign n2078 = ~n2076 & ~n2077;
  assign n2079 = 171 & 494;
  assign n2080 = ~n2078 & ~n2079;
  assign n2081 = ~n2078 & ~n2080;
  assign n2082 = ~n2079 & ~n2080;
  assign n2083 = ~n2081 & ~n2082;
  assign n2084 = ~n1994 & ~n1999;
  assign n2085 = ~n2083 & ~n2084;
  assign n2086 = ~n2083 & ~n2085;
  assign n2087 = ~n2084 & ~n2085;
  assign n2088 = ~n2086 & ~n2087;
  assign n2089 = 154 & 511;
  assign n2090 = ~n2088 & ~n2089;
  assign n2091 = ~n2088 & ~n2090;
  assign n2092 = ~n2089 & ~n2090;
  assign n2093 = ~n2091 & ~n2092;
  assign n2094 = ~n2004 & ~n2009;
  assign n2095 = ~n2093 & ~n2094;
  assign n2096 = ~n2093 & ~n2095;
  assign n2097 = ~n2094 & ~n2095;
  assign n2098 = ~n2096 & ~n2097;
  assign n2099 = 137 & 528;
  assign n2100 = ~n2098 & ~n2099;
  assign n2101 = ~n2098 & ~n2100;
  assign n2102 = ~n2099 & ~n2100;
  assign n2103 = ~n2101 & ~n2102;
  assign n2104 = ~n2014 & ~n2019;
  assign n2105 = ~n2103 & ~n2104;
  assign n2106 = ~n2103 & ~n2105;
  assign n2107 = ~n2104 & ~n2105;
  assign n2108 = ~n2106 & ~n2107;
  assign n2109 = ~n2024 & ~n2029;
  assign n2110 = ~n2108 & ~n2109;
  assign n2111 = ~n2108 & ~n2110;
  assign n2112 = ~n2109 & ~n2110;
  assign 6220 = ~n2111 & ~n2112;
  assign n2114 = 256 & 426;
  assign n2115 = ~n2035 & ~n2040;
  assign n2116 = ~n2114 & ~n2115;
  assign n2117 = ~n2114 & ~n2116;
  assign n2118 = ~n2115 & ~n2116;
  assign n2119 = ~n2117 & ~n2118;
  assign n2120 = 239 & 443;
  assign n2121 = ~n2119 & ~n2120;
  assign n2122 = ~n2119 & ~n2121;
  assign n2123 = ~n2120 & ~n2121;
  assign n2124 = ~n2122 & ~n2123;
  assign n2125 = ~n2045 & ~n2050;
  assign n2126 = ~n2124 & ~n2125;
  assign n2127 = ~n2124 & ~n2126;
  assign n2128 = ~n2125 & ~n2126;
  assign n2129 = ~n2127 & ~n2128;
  assign n2130 = 222 & 460;
  assign n2131 = ~n2129 & ~n2130;
  assign n2132 = ~n2129 & ~n2131;
  assign n2133 = ~n2130 & ~n2131;
  assign n2134 = ~n2132 & ~n2133;
  assign n2135 = ~n2055 & ~n2060;
  assign n2136 = ~n2134 & ~n2135;
  assign n2137 = ~n2134 & ~n2136;
  assign n2138 = ~n2135 & ~n2136;
  assign n2139 = ~n2137 & ~n2138;
  assign n2140 = 205 & 477;
  assign n2141 = ~n2139 & ~n2140;
  assign n2142 = ~n2139 & ~n2141;
  assign n2143 = ~n2140 & ~n2141;
  assign n2144 = ~n2142 & ~n2143;
  assign n2145 = ~n2065 & ~n2070;
  assign n2146 = ~n2144 & ~n2145;
  assign n2147 = ~n2144 & ~n2146;
  assign n2148 = ~n2145 & ~n2146;
  assign n2149 = ~n2147 & ~n2148;
  assign n2150 = 188 & 494;
  assign n2151 = ~n2149 & ~n2150;
  assign n2152 = ~n2149 & ~n2151;
  assign n2153 = ~n2150 & ~n2151;
  assign n2154 = ~n2152 & ~n2153;
  assign n2155 = ~n2075 & ~n2080;
  assign n2156 = ~n2154 & ~n2155;
  assign n2157 = ~n2154 & ~n2156;
  assign n2158 = ~n2155 & ~n2156;
  assign n2159 = ~n2157 & ~n2158;
  assign n2160 = 171 & 511;
  assign n2161 = ~n2159 & ~n2160;
  assign n2162 = ~n2159 & ~n2161;
  assign n2163 = ~n2160 & ~n2161;
  assign n2164 = ~n2162 & ~n2163;
  assign n2165 = ~n2085 & ~n2090;
  assign n2166 = ~n2164 & ~n2165;
  assign n2167 = ~n2164 & ~n2166;
  assign n2168 = ~n2165 & ~n2166;
  assign n2169 = ~n2167 & ~n2168;
  assign n2170 = 154 & 528;
  assign n2171 = ~n2169 & ~n2170;
  assign n2172 = ~n2169 & ~n2171;
  assign n2173 = ~n2170 & ~n2171;
  assign n2174 = ~n2172 & ~n2173;
  assign n2175 = ~n2095 & ~n2100;
  assign n2176 = ~n2174 & ~n2175;
  assign n2177 = ~n2174 & ~n2176;
  assign n2178 = ~n2175 & ~n2176;
  assign n2179 = ~n2177 & ~n2178;
  assign n2180 = ~n2105 & ~n2110;
  assign n2181 = ~n2179 & ~n2180;
  assign n2182 = ~n2179 & ~n2181;
  assign n2183 = ~n2180 & ~n2181;
  assign 6230 = ~n2182 & ~n2183;
  assign n2185 = 256 & 443;
  assign n2186 = ~n2116 & ~n2121;
  assign n2187 = ~n2185 & ~n2186;
  assign n2188 = ~n2185 & ~n2187;
  assign n2189 = ~n2186 & ~n2187;
  assign n2190 = ~n2188 & ~n2189;
  assign n2191 = 239 & 460;
  assign n2192 = ~n2190 & ~n2191;
  assign n2193 = ~n2190 & ~n2192;
  assign n2194 = ~n2191 & ~n2192;
  assign n2195 = ~n2193 & ~n2194;
  assign n2196 = ~n2126 & ~n2131;
  assign n2197 = ~n2195 & ~n2196;
  assign n2198 = ~n2195 & ~n2197;
  assign n2199 = ~n2196 & ~n2197;
  assign n2200 = ~n2198 & ~n2199;
  assign n2201 = 222 & 477;
  assign n2202 = ~n2200 & ~n2201;
  assign n2203 = ~n2200 & ~n2202;
  assign n2204 = ~n2201 & ~n2202;
  assign n2205 = ~n2203 & ~n2204;
  assign n2206 = ~n2136 & ~n2141;
  assign n2207 = ~n2205 & ~n2206;
  assign n2208 = ~n2205 & ~n2207;
  assign n2209 = ~n2206 & ~n2207;
  assign n2210 = ~n2208 & ~n2209;
  assign n2211 = 205 & 494;
  assign n2212 = ~n2210 & ~n2211;
  assign n2213 = ~n2210 & ~n2212;
  assign n2214 = ~n2211 & ~n2212;
  assign n2215 = ~n2213 & ~n2214;
  assign n2216 = ~n2146 & ~n2151;
  assign n2217 = ~n2215 & ~n2216;
  assign n2218 = ~n2215 & ~n2217;
  assign n2219 = ~n2216 & ~n2217;
  assign n2220 = ~n2218 & ~n2219;
  assign n2221 = 188 & 511;
  assign n2222 = ~n2220 & ~n2221;
  assign n2223 = ~n2220 & ~n2222;
  assign n2224 = ~n2221 & ~n2222;
  assign n2225 = ~n2223 & ~n2224;
  assign n2226 = ~n2156 & ~n2161;
  assign n2227 = ~n2225 & ~n2226;
  assign n2228 = ~n2225 & ~n2227;
  assign n2229 = ~n2226 & ~n2227;
  assign n2230 = ~n2228 & ~n2229;
  assign n2231 = 171 & 528;
  assign n2232 = ~n2230 & ~n2231;
  assign n2233 = ~n2230 & ~n2232;
  assign n2234 = ~n2231 & ~n2232;
  assign n2235 = ~n2233 & ~n2234;
  assign n2236 = ~n2166 & ~n2171;
  assign n2237 = ~n2235 & ~n2236;
  assign n2238 = ~n2235 & ~n2237;
  assign n2239 = ~n2236 & ~n2237;
  assign n2240 = ~n2238 & ~n2239;
  assign n2241 = ~n2176 & ~n2181;
  assign n2242 = ~n2240 & ~n2241;
  assign n2243 = ~n2240 & ~n2242;
  assign n2244 = ~n2241 & ~n2242;
  assign 6240 = ~n2243 & ~n2244;
  assign n2246 = 256 & 460;
  assign n2247 = ~n2187 & ~n2192;
  assign n2248 = ~n2246 & ~n2247;
  assign n2249 = ~n2246 & ~n2248;
  assign n2250 = ~n2247 & ~n2248;
  assign n2251 = ~n2249 & ~n2250;
  assign n2252 = 239 & 477;
  assign n2253 = ~n2251 & ~n2252;
  assign n2254 = ~n2251 & ~n2253;
  assign n2255 = ~n2252 & ~n2253;
  assign n2256 = ~n2254 & ~n2255;
  assign n2257 = ~n2197 & ~n2202;
  assign n2258 = ~n2256 & ~n2257;
  assign n2259 = ~n2256 & ~n2258;
  assign n2260 = ~n2257 & ~n2258;
  assign n2261 = ~n2259 & ~n2260;
  assign n2262 = 222 & 494;
  assign n2263 = ~n2261 & ~n2262;
  assign n2264 = ~n2261 & ~n2263;
  assign n2265 = ~n2262 & ~n2263;
  assign n2266 = ~n2264 & ~n2265;
  assign n2267 = ~n2207 & ~n2212;
  assign n2268 = ~n2266 & ~n2267;
  assign n2269 = ~n2266 & ~n2268;
  assign n2270 = ~n2267 & ~n2268;
  assign n2271 = ~n2269 & ~n2270;
  assign n2272 = 205 & 511;
  assign n2273 = ~n2271 & ~n2272;
  assign n2274 = ~n2271 & ~n2273;
  assign n2275 = ~n2272 & ~n2273;
  assign n2276 = ~n2274 & ~n2275;
  assign n2277 = ~n2217 & ~n2222;
  assign n2278 = ~n2276 & ~n2277;
  assign n2279 = ~n2276 & ~n2278;
  assign n2280 = ~n2277 & ~n2278;
  assign n2281 = ~n2279 & ~n2280;
  assign n2282 = 188 & 528;
  assign n2283 = ~n2281 & ~n2282;
  assign n2284 = ~n2281 & ~n2283;
  assign n2285 = ~n2282 & ~n2283;
  assign n2286 = ~n2284 & ~n2285;
  assign n2287 = ~n2227 & ~n2232;
  assign n2288 = ~n2286 & ~n2287;
  assign n2289 = ~n2286 & ~n2288;
  assign n2290 = ~n2287 & ~n2288;
  assign n2291 = ~n2289 & ~n2290;
  assign n2292 = ~n2237 & ~n2242;
  assign n2293 = ~n2291 & ~n2292;
  assign n2294 = ~n2291 & ~n2293;
  assign n2295 = ~n2292 & ~n2293;
  assign 6250 = ~n2294 & ~n2295;
  assign n2297 = 256 & 477;
  assign n2298 = ~n2248 & ~n2253;
  assign n2299 = ~n2297 & ~n2298;
  assign n2300 = ~n2297 & ~n2299;
  assign n2301 = ~n2298 & ~n2299;
  assign n2302 = ~n2300 & ~n2301;
  assign n2303 = 239 & 494;
  assign n2304 = ~n2302 & ~n2303;
  assign n2305 = ~n2302 & ~n2304;
  assign n2306 = ~n2303 & ~n2304;
  assign n2307 = ~n2305 & ~n2306;
  assign n2308 = ~n2258 & ~n2263;
  assign n2309 = ~n2307 & ~n2308;
  assign n2310 = ~n2307 & ~n2309;
  assign n2311 = ~n2308 & ~n2309;
  assign n2312 = ~n2310 & ~n2311;
  assign n2313 = 222 & 511;
  assign n2314 = ~n2312 & ~n2313;
  assign n2315 = ~n2312 & ~n2314;
  assign n2316 = ~n2313 & ~n2314;
  assign n2317 = ~n2315 & ~n2316;
  assign n2318 = ~n2268 & ~n2273;
  assign n2319 = ~n2317 & ~n2318;
  assign n2320 = ~n2317 & ~n2319;
  assign n2321 = ~n2318 & ~n2319;
  assign n2322 = ~n2320 & ~n2321;
  assign n2323 = 205 & 528;
  assign n2324 = ~n2322 & ~n2323;
  assign n2325 = ~n2322 & ~n2324;
  assign n2326 = ~n2323 & ~n2324;
  assign n2327 = ~n2325 & ~n2326;
  assign n2328 = ~n2278 & ~n2283;
  assign n2329 = ~n2327 & ~n2328;
  assign n2330 = ~n2327 & ~n2329;
  assign n2331 = ~n2328 & ~n2329;
  assign n2332 = ~n2330 & ~n2331;
  assign n2333 = ~n2288 & ~n2293;
  assign n2334 = ~n2332 & ~n2333;
  assign n2335 = ~n2332 & ~n2334;
  assign n2336 = ~n2333 & ~n2334;
  assign 6260 = ~n2335 & ~n2336;
  assign n2338 = 256 & 494;
  assign n2339 = ~n2299 & ~n2304;
  assign n2340 = ~n2338 & ~n2339;
  assign n2341 = ~n2338 & ~n2340;
  assign n2342 = ~n2339 & ~n2340;
  assign n2343 = ~n2341 & ~n2342;
  assign n2344 = 239 & 511;
  assign n2345 = ~n2343 & ~n2344;
  assign n2346 = ~n2343 & ~n2345;
  assign n2347 = ~n2344 & ~n2345;
  assign n2348 = ~n2346 & ~n2347;
  assign n2349 = ~n2309 & ~n2314;
  assign n2350 = ~n2348 & ~n2349;
  assign n2351 = ~n2348 & ~n2350;
  assign n2352 = ~n2349 & ~n2350;
  assign n2353 = ~n2351 & ~n2352;
  assign n2354 = 222 & 528;
  assign n2355 = ~n2353 & ~n2354;
  assign n2356 = ~n2353 & ~n2355;
  assign n2357 = ~n2354 & ~n2355;
  assign n2358 = ~n2356 & ~n2357;
  assign n2359 = ~n2319 & ~n2324;
  assign n2360 = ~n2358 & ~n2359;
  assign n2361 = ~n2358 & ~n2360;
  assign n2362 = ~n2359 & ~n2360;
  assign n2363 = ~n2361 & ~n2362;
  assign n2364 = ~n2329 & ~n2334;
  assign n2365 = ~n2363 & ~n2364;
  assign n2366 = ~n2363 & ~n2365;
  assign n2367 = ~n2364 & ~n2365;
  assign 6270 = ~n2366 & ~n2367;
  assign n2369 = 256 & 511;
  assign n2370 = ~n2340 & ~n2345;
  assign n2371 = ~n2369 & ~n2370;
  assign n2372 = ~n2369 & ~n2371;
  assign n2373 = ~n2370 & ~n2371;
  assign n2374 = ~n2372 & ~n2373;
  assign n2375 = 239 & 528;
  assign n2376 = ~n2374 & ~n2375;
  assign n2377 = ~n2374 & ~n2376;
  assign n2378 = ~n2375 & ~n2376;
  assign n2379 = ~n2377 & ~n2378;
  assign n2380 = ~n2350 & ~n2355;
  assign n2381 = ~n2379 & ~n2380;
  assign n2382 = ~n2379 & ~n2381;
  assign n2383 = ~n2380 & ~n2381;
  assign n2384 = ~n2382 & ~n2383;
  assign n2385 = ~n2360 & ~n2365;
  assign n2386 = ~n2384 & ~n2385;
  assign n2387 = ~n2384 & ~n2386;
  assign n2388 = ~n2385 & ~n2386;
  assign 6280 = ~n2387 & ~n2388;
  assign n2390 = 256 & 528;
  assign n2391 = ~n2371 & ~n2376;
  assign n2392 = ~n2390 & ~n2391;
  assign n2393 = ~n2390 & ~n2392;
  assign n2394 = ~n2391 & ~n2392;
  assign n2395 = ~n2393 & ~n2394;
  assign n2396 = ~n2381 & ~n2386;
  assign n2397 = ~n2395 & ~n2396;
  assign 6287 = ~n2392 & ~n2397;
  assign n2399 = ~n2395 & ~n2397;
  assign n2400 = ~n2396 & ~n2397;
  assign 6288 = ~n2399 & ~n2400;
endmodule
