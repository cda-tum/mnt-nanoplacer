module top (
    \in00 , \in01 , \in02 , \in03 , \in04 , \in05 , \in06 ,
    \in07 , \in08 , \in09 , \in010 , \in011 , \in012 ,
    \in013 , \in014 , \in015 , \in016 , \in017 , \in018 ,
    \in019 , \in020 , \in021 , \in022 , \in023 , \in024 ,
    \in025 , \in026 , \in027 , \in028 , \in029 , \in030 ,
    \in031 , \in032 , \in033 , \in034 , \in035 , \in036 ,
    \in037 , \in038 , \in039 , \in040 , \in041 , \in042 ,
    \in043 , \in044 , \in045 , \in046 , \in047 , \in048 ,
    \in049 , \in050 , \in051 , \in052 , \in053 , \in054 ,
    \in055 , \in056 , \in057 , \in058 , \in059 , \in060 ,
    \in061 , \in062 , \in063 , \in064 , \in065 , \in066 ,
    \in067 , \in068 , \in069 , \in070 , \in071 , \in072 ,
    \in073 , \in074 , \in075 , \in076 , \in077 , \in078 ,
    \in079 , \in080 , \in081 , \in082 , \in083 , \in084 ,
    \in085 , \in086 , \in087 , \in088 , \in089 , \in090 ,
    \in091 , \in092 , \in093 , \in094 , \in095 , \in096 ,
    \in097 , \in098 , \in099 , \in0100 , \in0101 , \in0102 ,
    \in0103 , \in0104 , \in0105 , \in0106 , \in0107 , \in0108 ,
    \in0109 , \in0110 , \in0111 , \in0112 , \in0113 , \in0114 ,
    \in0115 , \in0116 , \in0117 , \in0118 , \in0119 , \in0120 ,
    \in0121 , \in0122 , \in0123 , \in0124 , \in0125 , \in0126 ,
    \in0127 , \in10 , \in11 , \in12 , \in13 , \in14 , \in15 ,
    \in16 , \in17 , \in18 , \in19 , \in110 , \in111 ,
    \in112 , \in113 , \in114 , \in115 , \in116 , \in117 ,
    \in118 , \in119 , \in120 , \in121 , \in122 , \in123 ,
    \in124 , \in125 , \in126 , \in127 , \in128 , \in129 ,
    \in130 , \in131 , \in132 , \in133 , \in134 , \in135 ,
    \in136 , \in137 , \in138 , \in139 , \in140 , \in141 ,
    \in142 , \in143 , \in144 , \in145 , \in146 , \in147 ,
    \in148 , \in149 , \in150 , \in151 , \in152 , \in153 ,
    \in154 , \in155 , \in156 , \in157 , \in158 , \in159 ,
    \in160 , \in161 , \in162 , \in163 , \in164 , \in165 ,
    \in166 , \in167 , \in168 , \in169 , \in170 , \in171 ,
    \in172 , \in173 , \in174 , \in175 , \in176 , \in177 ,
    \in178 , \in179 , \in180 , \in181 , \in182 , \in183 ,
    \in184 , \in185 , \in186 , \in187 , \in188 , \in189 ,
    \in190 , \in191 , \in192 , \in193 , \in194 , \in195 ,
    \in196 , \in197 , \in198 , \in199 , \in1100 , \in1101 ,
    \in1102 , \in1103 , \in1104 , \in1105 , \in1106 , \in1107 ,
    \in1108 , \in1109 , \in1110 , \in1111 , \in1112 , \in1113 ,
    \in1114 , \in1115 , \in1116 , \in1117 , \in1118 , \in1119 ,
    \in1120 , \in1121 , \in1122 , \in1123 , \in1124 , \in1125 ,
    \in1126 , \in1127 , \in20 , \in21 , \in22 , \in23 ,
    \in24 , \in25 , \in26 , \in27 , \in28 , \in29 , \in210 ,
    \in211 , \in212 , \in213 , \in214 , \in215 , \in216 ,
    \in217 , \in218 , \in219 , \in220 , \in221 , \in222 ,
    \in223 , \in224 , \in225 , \in226 , \in227 , \in228 ,
    \in229 , \in230 , \in231 , \in232 , \in233 , \in234 ,
    \in235 , \in236 , \in237 , \in238 , \in239 , \in240 ,
    \in241 , \in242 , \in243 , \in244 , \in245 , \in246 ,
    \in247 , \in248 , \in249 , \in250 , \in251 , \in252 ,
    \in253 , \in254 , \in255 , \in256 , \in257 , \in258 ,
    \in259 , \in260 , \in261 , \in262 , \in263 , \in264 ,
    \in265 , \in266 , \in267 , \in268 , \in269 , \in270 ,
    \in271 , \in272 , \in273 , \in274 , \in275 , \in276 ,
    \in277 , \in278 , \in279 , \in280 , \in281 , \in282 ,
    \in283 , \in284 , \in285 , \in286 , \in287 , \in288 ,
    \in289 , \in290 , \in291 , \in292 , \in293 , \in294 ,
    \in295 , \in296 , \in297 , \in298 , \in299 , \in2100 ,
    \in2101 , \in2102 , \in2103 , \in2104 , \in2105 , \in2106 ,
    \in2107 , \in2108 , \in2109 , \in2110 , \in2111 , \in2112 ,
    \in2113 , \in2114 , \in2115 , \in2116 , \in2117 , \in2118 ,
    \in2119 , \in2120 , \in2121 , \in2122 , \in2123 , \in2124 ,
    \in2125 , \in2126 , \in2127 , \in30 , \in31 , \in32 ,
    \in33 , \in34 , \in35 , \in36 , \in37 , \in38 , \in39 ,
    \in310 , \in311 , \in312 , \in313 , \in314 , \in315 ,
    \in316 , \in317 , \in318 , \in319 , \in320 , \in321 ,
    \in322 , \in323 , \in324 , \in325 , \in326 , \in327 ,
    \in328 , \in329 , \in330 , \in331 , \in332 , \in333 ,
    \in334 , \in335 , \in336 , \in337 , \in338 , \in339 ,
    \in340 , \in341 , \in342 , \in343 , \in344 , \in345 ,
    \in346 , \in347 , \in348 , \in349 , \in350 , \in351 ,
    \in352 , \in353 , \in354 , \in355 , \in356 , \in357 ,
    \in358 , \in359 , \in360 , \in361 , \in362 , \in363 ,
    \in364 , \in365 , \in366 , \in367 , \in368 , \in369 ,
    \in370 , \in371 , \in372 , \in373 , \in374 , \in375 ,
    \in376 , \in377 , \in378 , \in379 , \in380 , \in381 ,
    \in382 , \in383 , \in384 , \in385 , \in386 , \in387 ,
    \in388 , \in389 , \in390 , \in391 , \in392 , \in393 ,
    \in394 , \in395 , \in396 , \in397 , \in398 , \in399 ,
    \in3100 , \in3101 , \in3102 , \in3103 , \in3104 , \in3105 ,
    \in3106 , \in3107 , \in3108 , \in3109 , \in3110 , \in3111 ,
    \in3112 , \in3113 , \in3114 , \in3115 , \in3116 , \in3117 ,
    \in3118 , \in3119 , \in3120 , \in3121 , \in3122 , \in3123 ,
    \in3124 , \in3125 , \in3126 , \in3127 ,
    \result0 , \result1 , \result2 , \result3 , \result4 ,
    \result5 , \result6 , \result7 , \result8 , \result9 ,
    \result10 , \result11 , \result12 , \result13 , \result14 ,
    \result15 , \result16 , \result17 , \result18 , \result19 ,
    \result20 , \result21 , \result22 , \result23 , \result24 ,
    \result25 , \result26 , \result27 , \result28 , \result29 ,
    \result30 , \result31 , \result32 , \result33 , \result34 ,
    \result35 , \result36 , \result37 , \result38 , \result39 ,
    \result40 , \result41 , \result42 , \result43 , \result44 ,
    \result45 , \result46 , \result47 , \result48 , \result49 ,
    \result50 , \result51 , \result52 , \result53 , \result54 ,
    \result55 , \result56 , \result57 , \result58 , \result59 ,
    \result60 , \result61 , \result62 , \result63 , \result64 ,
    \result65 , \result66 , \result67 , \result68 , \result69 ,
    \result70 , \result71 , \result72 , \result73 , \result74 ,
    \result75 , \result76 , \result77 , \result78 , \result79 ,
    \result80 , \result81 , \result82 , \result83 , \result84 ,
    \result85 , \result86 , \result87 , \result88 , \result89 ,
    \result90 , \result91 , \result92 , \result93 , \result94 ,
    \result95 , \result96 , \result97 , \result98 , \result99 ,
    \result100 , \result101 , \result102 , \result103 ,
    \result104 , \result105 , \result106 , \result107 ,
    \result108 , \result109 , \result110 , \result111 ,
    \result112 , \result113 , \result114 , \result115 ,
    \result116 , \result117 , \result118 , \result119 ,
    \result120 , \result121 , \result122 , \result123 ,
    \result124 , \result125 , \result126 , \result127 ,
    \address0 , \address1   );
  input  \in00 , \in01 , \in02 , \in03 , \in04 , \in05 ,
    \in06 , \in07 , \in08 , \in09 , \in010 , \in011 ,
    \in012 , \in013 , \in014 , \in015 , \in016 , \in017 ,
    \in018 , \in019 , \in020 , \in021 , \in022 , \in023 ,
    \in024 , \in025 , \in026 , \in027 , \in028 , \in029 ,
    \in030 , \in031 , \in032 , \in033 , \in034 , \in035 ,
    \in036 , \in037 , \in038 , \in039 , \in040 , \in041 ,
    \in042 , \in043 , \in044 , \in045 , \in046 , \in047 ,
    \in048 , \in049 , \in050 , \in051 , \in052 , \in053 ,
    \in054 , \in055 , \in056 , \in057 , \in058 , \in059 ,
    \in060 , \in061 , \in062 , \in063 , \in064 , \in065 ,
    \in066 , \in067 , \in068 , \in069 , \in070 , \in071 ,
    \in072 , \in073 , \in074 , \in075 , \in076 , \in077 ,
    \in078 , \in079 , \in080 , \in081 , \in082 , \in083 ,
    \in084 , \in085 , \in086 , \in087 , \in088 , \in089 ,
    \in090 , \in091 , \in092 , \in093 , \in094 , \in095 ,
    \in096 , \in097 , \in098 , \in099 , \in0100 , \in0101 ,
    \in0102 , \in0103 , \in0104 , \in0105 , \in0106 , \in0107 ,
    \in0108 , \in0109 , \in0110 , \in0111 , \in0112 , \in0113 ,
    \in0114 , \in0115 , \in0116 , \in0117 , \in0118 , \in0119 ,
    \in0120 , \in0121 , \in0122 , \in0123 , \in0124 , \in0125 ,
    \in0126 , \in0127 , \in10 , \in11 , \in12 , \in13 ,
    \in14 , \in15 , \in16 , \in17 , \in18 , \in19 , \in110 ,
    \in111 , \in112 , \in113 , \in114 , \in115 , \in116 ,
    \in117 , \in118 , \in119 , \in120 , \in121 , \in122 ,
    \in123 , \in124 , \in125 , \in126 , \in127 , \in128 ,
    \in129 , \in130 , \in131 , \in132 , \in133 , \in134 ,
    \in135 , \in136 , \in137 , \in138 , \in139 , \in140 ,
    \in141 , \in142 , \in143 , \in144 , \in145 , \in146 ,
    \in147 , \in148 , \in149 , \in150 , \in151 , \in152 ,
    \in153 , \in154 , \in155 , \in156 , \in157 , \in158 ,
    \in159 , \in160 , \in161 , \in162 , \in163 , \in164 ,
    \in165 , \in166 , \in167 , \in168 , \in169 , \in170 ,
    \in171 , \in172 , \in173 , \in174 , \in175 , \in176 ,
    \in177 , \in178 , \in179 , \in180 , \in181 , \in182 ,
    \in183 , \in184 , \in185 , \in186 , \in187 , \in188 ,
    \in189 , \in190 , \in191 , \in192 , \in193 , \in194 ,
    \in195 , \in196 , \in197 , \in198 , \in199 , \in1100 ,
    \in1101 , \in1102 , \in1103 , \in1104 , \in1105 , \in1106 ,
    \in1107 , \in1108 , \in1109 , \in1110 , \in1111 , \in1112 ,
    \in1113 , \in1114 , \in1115 , \in1116 , \in1117 , \in1118 ,
    \in1119 , \in1120 , \in1121 , \in1122 , \in1123 , \in1124 ,
    \in1125 , \in1126 , \in1127 , \in20 , \in21 , \in22 ,
    \in23 , \in24 , \in25 , \in26 , \in27 , \in28 , \in29 ,
    \in210 , \in211 , \in212 , \in213 , \in214 , \in215 ,
    \in216 , \in217 , \in218 , \in219 , \in220 , \in221 ,
    \in222 , \in223 , \in224 , \in225 , \in226 , \in227 ,
    \in228 , \in229 , \in230 , \in231 , \in232 , \in233 ,
    \in234 , \in235 , \in236 , \in237 , \in238 , \in239 ,
    \in240 , \in241 , \in242 , \in243 , \in244 , \in245 ,
    \in246 , \in247 , \in248 , \in249 , \in250 , \in251 ,
    \in252 , \in253 , \in254 , \in255 , \in256 , \in257 ,
    \in258 , \in259 , \in260 , \in261 , \in262 , \in263 ,
    \in264 , \in265 , \in266 , \in267 , \in268 , \in269 ,
    \in270 , \in271 , \in272 , \in273 , \in274 , \in275 ,
    \in276 , \in277 , \in278 , \in279 , \in280 , \in281 ,
    \in282 , \in283 , \in284 , \in285 , \in286 , \in287 ,
    \in288 , \in289 , \in290 , \in291 , \in292 , \in293 ,
    \in294 , \in295 , \in296 , \in297 , \in298 , \in299 ,
    \in2100 , \in2101 , \in2102 , \in2103 , \in2104 , \in2105 ,
    \in2106 , \in2107 , \in2108 , \in2109 , \in2110 , \in2111 ,
    \in2112 , \in2113 , \in2114 , \in2115 , \in2116 , \in2117 ,
    \in2118 , \in2119 , \in2120 , \in2121 , \in2122 , \in2123 ,
    \in2124 , \in2125 , \in2126 , \in2127 , \in30 , \in31 ,
    \in32 , \in33 , \in34 , \in35 , \in36 , \in37 , \in38 ,
    \in39 , \in310 , \in311 , \in312 , \in313 , \in314 ,
    \in315 , \in316 , \in317 , \in318 , \in319 , \in320 ,
    \in321 , \in322 , \in323 , \in324 , \in325 , \in326 ,
    \in327 , \in328 , \in329 , \in330 , \in331 , \in332 ,
    \in333 , \in334 , \in335 , \in336 , \in337 , \in338 ,
    \in339 , \in340 , \in341 , \in342 , \in343 , \in344 ,
    \in345 , \in346 , \in347 , \in348 , \in349 , \in350 ,
    \in351 , \in352 , \in353 , \in354 , \in355 , \in356 ,
    \in357 , \in358 , \in359 , \in360 , \in361 , \in362 ,
    \in363 , \in364 , \in365 , \in366 , \in367 , \in368 ,
    \in369 , \in370 , \in371 , \in372 , \in373 , \in374 ,
    \in375 , \in376 , \in377 , \in378 , \in379 , \in380 ,
    \in381 , \in382 , \in383 , \in384 , \in385 , \in386 ,
    \in387 , \in388 , \in389 , \in390 , \in391 , \in392 ,
    \in393 , \in394 , \in395 , \in396 , \in397 , \in398 ,
    \in399 , \in3100 , \in3101 , \in3102 , \in3103 , \in3104 ,
    \in3105 , \in3106 , \in3107 , \in3108 , \in3109 , \in3110 ,
    \in3111 , \in3112 , \in3113 , \in3114 , \in3115 , \in3116 ,
    \in3117 , \in3118 , \in3119 , \in3120 , \in3121 , \in3122 ,
    \in3123 , \in3124 , \in3125 , \in3126 , \in3127 ;
  output \result0 , \result1 , \result2 , \result3 , \result4 ,
    \result5 , \result6 , \result7 , \result8 , \result9 ,
    \result10 , \result11 , \result12 , \result13 , \result14 ,
    \result15 , \result16 , \result17 , \result18 , \result19 ,
    \result20 , \result21 , \result22 , \result23 , \result24 ,
    \result25 , \result26 , \result27 , \result28 , \result29 ,
    \result30 , \result31 , \result32 , \result33 , \result34 ,
    \result35 , \result36 , \result37 , \result38 , \result39 ,
    \result40 , \result41 , \result42 , \result43 , \result44 ,
    \result45 , \result46 , \result47 , \result48 , \result49 ,
    \result50 , \result51 , \result52 , \result53 , \result54 ,
    \result55 , \result56 , \result57 , \result58 , \result59 ,
    \result60 , \result61 , \result62 , \result63 , \result64 ,
    \result65 , \result66 , \result67 , \result68 , \result69 ,
    \result70 , \result71 , \result72 , \result73 , \result74 ,
    \result75 , \result76 , \result77 , \result78 , \result79 ,
    \result80 , \result81 , \result82 , \result83 , \result84 ,
    \result85 , \result86 , \result87 , \result88 , \result89 ,
    \result90 , \result91 , \result92 , \result93 , \result94 ,
    \result95 , \result96 , \result97 , \result98 , \result99 ,
    \result100 , \result101 , \result102 , \result103 ,
    \result104 , \result105 , \result106 , \result107 ,
    \result108 , \result109 , \result110 , \result111 ,
    \result112 , \result113 , \result114 , \result115 ,
    \result116 , \result117 , \result118 , \result119 ,
    \result120 , \result121 , \result122 , \result123 ,
    \result124 , \result125 , \result126 , \result127 ,
    \address0 , \address1 ;
  wire n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
    n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
    n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
    n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
    n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
    n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
    n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
    n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
    n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
    n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
    n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
    n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
    n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797,
    n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809,
    n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821,
    n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
    n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845,
    n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857,
    n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869,
    n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
    n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
    n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
    n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
    n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929,
    n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941,
    n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953,
    n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965,
    n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977,
    n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989,
    n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000,
    n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
    n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020,
    n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030,
    n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040,
    n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050,
    n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060,
    n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070,
    n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080,
    n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090,
    n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100,
    n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110,
    n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120,
    n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130,
    n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140,
    n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150,
    n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160,
    n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170,
    n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180,
    n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190,
    n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200,
    n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210,
    n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220,
    n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230,
    n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240,
    n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250,
    n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260,
    n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270,
    n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280,
    n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290,
    n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300,
    n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310,
    n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320,
    n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330,
    n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340,
    n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350,
    n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360,
    n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370,
    n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380,
    n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390,
    n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400,
    n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410,
    n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420,
    n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430,
    n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440,
    n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450,
    n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460,
    n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470,
    n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480,
    n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490,
    n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500,
    n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510,
    n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520,
    n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530,
    n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540,
    n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550,
    n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560,
    n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570,
    n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580,
    n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590,
    n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600,
    n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610,
    n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620,
    n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630,
    n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640,
    n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650,
    n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660,
    n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670,
    n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680,
    n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690,
    n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700,
    n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710,
    n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720,
    n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730,
    n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740,
    n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750,
    n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760,
    n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770,
    n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780,
    n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790,
    n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800,
    n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810,
    n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820,
    n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830,
    n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840,
    n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850,
    n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860,
    n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870,
    n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880,
    n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890,
    n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900,
    n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910,
    n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920,
    n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930,
    n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940,
    n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950,
    n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960,
    n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970,
    n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980,
    n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990,
    n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000,
    n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010,
    n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020,
    n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030,
    n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040,
    n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050,
    n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060,
    n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070,
    n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080,
    n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090,
    n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100,
    n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110,
    n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120,
    n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130,
    n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140,
    n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150,
    n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160,
    n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170,
    n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180,
    n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190,
    n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200,
    n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210,
    n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220,
    n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230,
    n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240,
    n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250,
    n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260,
    n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270,
    n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280,
    n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290,
    n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300,
    n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310,
    n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320,
    n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330,
    n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340,
    n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350,
    n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360,
    n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370,
    n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380,
    n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390,
    n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400,
    n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410,
    n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420,
    n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430,
    n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440,
    n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450,
    n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460,
    n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470,
    n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480,
    n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490,
    n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500,
    n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510,
    n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520,
    n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530,
    n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540,
    n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550,
    n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560,
    n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570,
    n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580,
    n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590,
    n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600,
    n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610,
    n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620,
    n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630,
    n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640,
    n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650,
    n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660,
    n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670,
    n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680,
    n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690,
    n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700,
    n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710,
    n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720,
    n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730,
    n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740,
    n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750,
    n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760,
    n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770,
    n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780,
    n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790,
    n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800,
    n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810,
    n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820,
    n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830,
    n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840,
    n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850,
    n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860,
    n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870,
    n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880,
    n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890,
    n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900,
    n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910,
    n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920,
    n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930,
    n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940,
    n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950,
    n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960,
    n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970,
    n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980,
    n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990,
    n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000,
    n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010,
    n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020,
    n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030,
    n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040,
    n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050,
    n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060,
    n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070,
    n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080,
    n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090,
    n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100,
    n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110,
    n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120,
    n3122, n3123, n3125, n3126, n3128, n3129, n3131, n3132, n3134, n3135,
    n3137, n3138, n3140, n3141, n3143, n3144, n3146, n3147, n3149, n3150,
    n3152, n3153, n3155, n3156, n3158, n3159, n3161, n3162, n3164, n3165,
    n3167, n3168, n3170, n3171, n3173, n3174, n3176, n3177, n3179, n3180,
    n3182, n3183, n3185, n3186, n3188, n3189, n3191, n3192, n3194, n3195,
    n3197, n3198, n3200, n3201, n3203, n3204, n3206, n3207, n3209, n3210,
    n3212, n3213, n3215, n3216, n3218, n3219, n3221, n3222, n3224, n3225,
    n3227, n3228, n3230, n3231, n3233, n3234, n3236, n3237, n3239, n3240,
    n3242, n3243, n3245, n3246, n3248, n3249, n3251, n3252, n3254, n3255,
    n3257, n3258, n3260, n3261, n3263, n3264, n3266, n3267, n3269, n3270,
    n3272, n3273, n3275, n3276, n3278, n3279, n3281, n3282, n3284, n3285,
    n3287, n3288, n3290, n3291, n3293, n3294, n3296, n3297, n3299, n3300,
    n3302, n3303, n3305, n3306, n3308, n3309, n3311, n3312, n3314, n3315,
    n3317, n3318, n3320, n3321, n3323, n3324, n3326, n3327, n3329, n3330,
    n3332, n3333, n3335, n3336, n3338, n3339, n3341, n3342, n3344, n3345,
    n3347, n3348, n3350, n3351, n3353, n3354, n3356, n3357, n3359, n3360,
    n3362, n3363, n3365, n3366, n3368, n3369, n3371, n3372, n3374, n3375,
    n3377, n3378, n3380, n3381, n3383, n3384, n3386, n3387, n3389, n3390,
    n3392, n3393, n3395, n3396, n3398, n3399, n3401, n3402, n3404, n3405,
    n3407, n3408, n3410, n3411, n3413, n3414, n3416, n3417, n3419, n3420,
    n3422, n3423, n3425, n3426, n3428, n3429, n3431, n3432, n3434, n3435,
    n3437, n3438, n3440, n3441, n3443, n3444, n3446, n3447, n3449, n3450,
    n3452, n3453, n3455, n3456, n3458, n3459, n3461, n3462, n3464, n3465,
    n3467, n3468, n3470, n3471, n3473, n3474, n3476, n3477, n3479, n3480,
    n3482, n3483, n3485, n3486, n3488, n3489, n3491, n3492, n3494, n3495,
    n3497, n3498, n3500, n3501, n3503, n3505, n3506;
  assign n643 = \in2119  & ~\in3119 ;
  assign n644 = ~\in2119  & \in3119 ;
  assign n645 = ~\in2118  & \in3118 ;
  assign n646 = ~n644 & ~n645;
  assign n647 = ~\in2117  & \in3117 ;
  assign n648 = \in2116  & ~\in3116 ;
  assign n649 = ~n647 & n648;
  assign n650 = \in2117  & ~\in3117 ;
  assign n651 = ~n649 & ~n650;
  assign n652 = n646 & ~n651;
  assign n653 = ~\in3118  & ~n644;
  assign n654 = \in2118  & n653;
  assign n655 = ~\in2112  & \in3112 ;
  assign n656 = ~\in2115  & \in3115 ;
  assign n657 = ~\in2114  & \in3114 ;
  assign n658 = ~n656 & ~n657;
  assign n659 = ~\in2113  & \in3113 ;
  assign n660 = \in2111  & ~\in3111 ;
  assign n661 = ~\in2111  & \in3111 ;
  assign n662 = ~\in2110  & \in3110 ;
  assign n663 = ~n661 & ~n662;
  assign n664 = ~\in2109  & \in3109 ;
  assign n665 = \in2108  & ~\in3108 ;
  assign n666 = ~n664 & n665;
  assign n667 = \in2109  & ~\in3109 ;
  assign n668 = ~n666 & ~n667;
  assign n669 = n663 & ~n668;
  assign n670 = ~\in3110  & ~n661;
  assign n671 = \in2110  & n670;
  assign n672 = \in2103  & ~\in3103 ;
  assign n673 = ~\in2103  & \in3103 ;
  assign n674 = ~\in2102  & \in3102 ;
  assign n675 = ~n673 & ~n674;
  assign n676 = ~\in2101  & \in3101 ;
  assign n677 = \in2100  & ~\in3100 ;
  assign n678 = ~n676 & n677;
  assign n679 = \in2101  & ~\in3101 ;
  assign n680 = ~n678 & ~n679;
  assign n681 = n675 & ~n680;
  assign n682 = ~\in3102  & ~n673;
  assign n683 = \in2102  & n682;
  assign n684 = ~\in296  & \in396 ;
  assign n685 = ~\in299  & \in399 ;
  assign n686 = ~\in298  & \in398 ;
  assign n687 = ~n685 & ~n686;
  assign n688 = ~\in297  & \in397 ;
  assign n689 = \in295  & ~\in395 ;
  assign n690 = ~\in295  & \in395 ;
  assign n691 = ~\in294  & \in394 ;
  assign n692 = ~n690 & ~n691;
  assign n693 = ~\in293  & \in393 ;
  assign n694 = \in292  & ~\in392 ;
  assign n695 = ~n693 & n694;
  assign n696 = \in293  & ~\in393 ;
  assign n697 = ~n695 & ~n696;
  assign n698 = n692 & ~n697;
  assign n699 = ~\in394  & ~n690;
  assign n700 = \in294  & n699;
  assign n701 = \in287  & ~\in387 ;
  assign n702 = ~\in287  & \in387 ;
  assign n703 = ~\in286  & \in386 ;
  assign n704 = ~n702 & ~n703;
  assign n705 = ~\in285  & \in385 ;
  assign n706 = \in284  & ~\in384 ;
  assign n707 = ~n705 & n706;
  assign n708 = \in285  & ~\in385 ;
  assign n709 = ~n707 & ~n708;
  assign n710 = n704 & ~n709;
  assign n711 = ~\in386  & ~n702;
  assign n712 = \in286  & n711;
  assign n713 = ~\in280  & \in380 ;
  assign n714 = ~\in283  & \in383 ;
  assign n715 = ~\in282  & \in382 ;
  assign n716 = ~n714 & ~n715;
  assign n717 = ~\in281  & \in381 ;
  assign n718 = \in279  & ~\in379 ;
  assign n719 = ~\in279  & \in379 ;
  assign n720 = ~\in278  & \in378 ;
  assign n721 = ~n719 & ~n720;
  assign n722 = ~\in277  & \in377 ;
  assign n723 = \in276  & ~\in376 ;
  assign n724 = ~n722 & n723;
  assign n725 = \in277  & ~\in377 ;
  assign n726 = ~n724 & ~n725;
  assign n727 = n721 & ~n726;
  assign n728 = ~\in378  & ~n719;
  assign n729 = \in278  & n728;
  assign n730 = \in271  & ~\in371 ;
  assign n731 = ~\in271  & \in371 ;
  assign n732 = ~\in270  & \in370 ;
  assign n733 = ~n731 & ~n732;
  assign n734 = ~\in269  & \in369 ;
  assign n735 = \in268  & ~\in368 ;
  assign n736 = ~n734 & n735;
  assign n737 = \in269  & ~\in369 ;
  assign n738 = ~n736 & ~n737;
  assign n739 = n733 & ~n738;
  assign n740 = ~\in370  & ~n731;
  assign n741 = \in270  & n740;
  assign n742 = ~\in267  & \in367 ;
  assign n743 = ~\in266  & \in366 ;
  assign n744 = ~n742 & ~n743;
  assign n745 = ~\in265  & \in365 ;
  assign n746 = \in263  & ~\in363 ;
  assign n747 = ~\in263  & \in363 ;
  assign n748 = ~\in262  & \in362 ;
  assign n749 = ~n747 & ~n748;
  assign n750 = ~\in260  & \in360 ;
  assign n751 = ~\in261  & \in361 ;
  assign n752 = ~n750 & ~n751;
  assign n753 = n749 & n752;
  assign n754 = \in259  & ~\in359 ;
  assign n755 = ~\in259  & \in359 ;
  assign n756 = ~\in258  & \in358 ;
  assign n757 = ~n755 & ~n756;
  assign n758 = ~\in257  & \in357 ;
  assign n759 = \in256  & ~\in356 ;
  assign n760 = ~n758 & n759;
  assign n761 = \in257  & ~\in357 ;
  assign n762 = ~n760 & ~n761;
  assign n763 = \in258  & ~\in358 ;
  assign n764 = n762 & ~n763;
  assign n765 = n757 & ~n764;
  assign n766 = ~n754 & ~n765;
  assign n767 = n753 & ~n766;
  assign n768 = \in260  & ~\in360 ;
  assign n769 = ~n751 & n768;
  assign n770 = \in261  & ~\in361 ;
  assign n771 = ~n769 & ~n770;
  assign n772 = n749 & ~n771;
  assign n773 = ~\in362  & ~n747;
  assign n774 = \in262  & n773;
  assign n775 = \in247  & ~\in347 ;
  assign n776 = ~\in247  & \in347 ;
  assign n777 = ~\in246  & \in346 ;
  assign n778 = ~n776 & ~n777;
  assign n779 = ~\in244  & \in344 ;
  assign n780 = ~\in245  & \in345 ;
  assign n781 = ~n779 & ~n780;
  assign n782 = n778 & n781;
  assign n783 = \in243  & ~\in343 ;
  assign n784 = ~\in243  & \in343 ;
  assign n785 = ~\in242  & \in342 ;
  assign n786 = ~n784 & ~n785;
  assign n787 = ~\in241  & \in341 ;
  assign n788 = \in240  & ~\in340 ;
  assign n789 = ~n787 & n788;
  assign n790 = \in241  & ~\in341 ;
  assign n791 = ~n789 & ~n790;
  assign n792 = \in242  & ~\in342 ;
  assign n793 = n791 & ~n792;
  assign n794 = n786 & ~n793;
  assign n795 = ~n783 & ~n794;
  assign n796 = n782 & ~n795;
  assign n797 = \in244  & ~\in344 ;
  assign n798 = ~n780 & n797;
  assign n799 = \in245  & ~\in345 ;
  assign n800 = ~n798 & ~n799;
  assign n801 = n778 & ~n800;
  assign n802 = ~\in346  & ~n776;
  assign n803 = \in246  & n802;
  assign n804 = ~\in232  & \in332 ;
  assign n805 = ~\in231  & \in331 ;
  assign n806 = ~\in230  & \in330 ;
  assign n807 = ~\in229  & \in329 ;
  assign n808 = ~\in228  & \in328 ;
  assign n809 = ~\in227  & \in327 ;
  assign n810 = ~\in226  & \in326 ;
  assign n811 = ~\in223  & \in323 ;
  assign n812 = ~\in222  & \in322 ;
  assign n813 = ~\in221  & \in321 ;
  assign n814 = ~\in220  & \in320 ;
  assign n815 = ~\in219  & \in319 ;
  assign n816 = ~\in218  & \in318 ;
  assign n817 = ~\in215  & \in315 ;
  assign n818 = ~\in214  & \in314 ;
  assign n819 = ~\in213  & \in313 ;
  assign n820 = ~\in212  & \in312 ;
  assign n821 = ~\in211  & \in311 ;
  assign n822 = ~\in210  & \in310 ;
  assign n823 = ~\in27  & \in37 ;
  assign n824 = ~\in26  & \in36 ;
  assign n825 = ~\in23  & \in33 ;
  assign n826 = \in20  & ~\in30 ;
  assign n827 = \in21  & n826;
  assign n828 = \in31  & ~n827;
  assign n829 = ~\in22  & \in32 ;
  assign n830 = ~\in21  & ~n826;
  assign n831 = ~n829 & ~n830;
  assign n832 = ~n828 & n831;
  assign n833 = \in22  & ~\in32 ;
  assign n834 = ~n832 & ~n833;
  assign n835 = ~n825 & ~n834;
  assign n836 = \in23  & ~\in33 ;
  assign n837 = ~n835 & ~n836;
  assign n838 = ~\in24  & n837;
  assign n839 = ~\in34  & ~n838;
  assign n840 = \in24  & ~n837;
  assign n841 = ~n839 & ~n840;
  assign n842 = ~\in25  & n841;
  assign n843 = ~\in35  & ~n842;
  assign n844 = \in25  & ~n841;
  assign n845 = ~n843 & ~n844;
  assign n846 = ~n824 & ~n845;
  assign n847 = \in26  & ~\in36 ;
  assign n848 = ~n846 & ~n847;
  assign n849 = ~n823 & ~n848;
  assign n850 = \in27  & ~\in37 ;
  assign n851 = ~n849 & ~n850;
  assign n852 = ~\in28  & n851;
  assign n853 = ~\in38  & ~n852;
  assign n854 = \in28  & ~n851;
  assign n855 = ~n853 & ~n854;
  assign n856 = ~\in29  & n855;
  assign n857 = ~\in39  & ~n856;
  assign n858 = \in29  & ~n855;
  assign n859 = ~n857 & ~n858;
  assign n860 = ~n822 & ~n859;
  assign n861 = \in210  & ~\in310 ;
  assign n862 = ~n860 & ~n861;
  assign n863 = ~n821 & ~n862;
  assign n864 = \in211  & ~\in311 ;
  assign n865 = ~n863 & ~n864;
  assign n866 = ~n820 & ~n865;
  assign n867 = \in212  & ~\in312 ;
  assign n868 = ~n866 & ~n867;
  assign n869 = ~n819 & ~n868;
  assign n870 = \in213  & ~\in313 ;
  assign n871 = ~n869 & ~n870;
  assign n872 = ~n818 & ~n871;
  assign n873 = \in214  & ~\in314 ;
  assign n874 = ~n872 & ~n873;
  assign n875 = ~n817 & ~n874;
  assign n876 = \in215  & ~\in315 ;
  assign n877 = ~n875 & ~n876;
  assign n878 = ~\in216  & n877;
  assign n879 = ~\in316  & ~n878;
  assign n880 = \in216  & ~n877;
  assign n881 = ~n879 & ~n880;
  assign n882 = ~\in217  & n881;
  assign n883 = ~\in317  & ~n882;
  assign n884 = \in217  & ~n881;
  assign n885 = ~n883 & ~n884;
  assign n886 = ~n816 & ~n885;
  assign n887 = \in218  & ~\in318 ;
  assign n888 = ~n886 & ~n887;
  assign n889 = ~n815 & ~n888;
  assign n890 = \in219  & ~\in319 ;
  assign n891 = ~n889 & ~n890;
  assign n892 = ~n814 & ~n891;
  assign n893 = \in220  & ~\in320 ;
  assign n894 = ~n892 & ~n893;
  assign n895 = ~n813 & ~n894;
  assign n896 = \in221  & ~\in321 ;
  assign n897 = ~n895 & ~n896;
  assign n898 = ~n812 & ~n897;
  assign n899 = \in222  & ~\in322 ;
  assign n900 = ~n898 & ~n899;
  assign n901 = ~n811 & ~n900;
  assign n902 = \in223  & ~\in323 ;
  assign n903 = ~n901 & ~n902;
  assign n904 = ~\in224  & n903;
  assign n905 = ~\in324  & ~n904;
  assign n906 = \in224  & ~n903;
  assign n907 = ~n905 & ~n906;
  assign n908 = ~\in225  & n907;
  assign n909 = ~\in325  & ~n908;
  assign n910 = \in225  & ~n907;
  assign n911 = ~n909 & ~n910;
  assign n912 = ~n810 & ~n911;
  assign n913 = \in226  & ~\in326 ;
  assign n914 = ~n912 & ~n913;
  assign n915 = ~n809 & ~n914;
  assign n916 = \in227  & ~\in327 ;
  assign n917 = ~n915 & ~n916;
  assign n918 = ~n808 & ~n917;
  assign n919 = \in228  & ~\in328 ;
  assign n920 = ~n918 & ~n919;
  assign n921 = ~n807 & ~n920;
  assign n922 = \in229  & ~\in329 ;
  assign n923 = ~n921 & ~n922;
  assign n924 = ~n806 & ~n923;
  assign n925 = \in230  & ~\in330 ;
  assign n926 = ~n924 & ~n925;
  assign n927 = ~n805 & ~n926;
  assign n928 = \in231  & ~\in331 ;
  assign n929 = ~n927 & ~n928;
  assign n930 = ~\in239  & \in339 ;
  assign n931 = ~\in238  & \in338 ;
  assign n932 = ~n930 & ~n931;
  assign n933 = ~\in236  & \in336 ;
  assign n934 = ~\in237  & \in337 ;
  assign n935 = ~n933 & ~n934;
  assign n936 = n932 & n935;
  assign n937 = ~\in233  & \in333 ;
  assign n938 = ~\in235  & \in335 ;
  assign n939 = ~\in234  & \in334 ;
  assign n940 = ~n938 & ~n939;
  assign n941 = ~n937 & n940;
  assign n942 = n936 & n941;
  assign n943 = ~n929 & n942;
  assign n944 = ~n804 & n943;
  assign n945 = \in239  & ~\in339 ;
  assign n946 = \in236  & ~\in336 ;
  assign n947 = ~n934 & n946;
  assign n948 = \in237  & ~\in337 ;
  assign n949 = ~n947 & ~n948;
  assign n950 = n932 & ~n949;
  assign n951 = ~\in338  & ~n930;
  assign n952 = \in238  & n951;
  assign n953 = \in235  & ~\in335 ;
  assign n954 = ~\in332  & ~n937;
  assign n955 = \in232  & n954;
  assign n956 = \in233  & ~\in333 ;
  assign n957 = ~n955 & ~n956;
  assign n958 = \in234  & ~\in334 ;
  assign n959 = n957 & ~n958;
  assign n960 = n940 & ~n959;
  assign n961 = ~n953 & ~n960;
  assign n962 = n936 & ~n961;
  assign n963 = ~n952 & ~n962;
  assign n964 = ~n950 & n963;
  assign n965 = ~n945 & n964;
  assign n966 = ~n944 & n965;
  assign n967 = ~\in240  & \in340 ;
  assign n968 = ~n787 & ~n967;
  assign n969 = n786 & n968;
  assign n970 = n782 & n969;
  assign n971 = ~n966 & n970;
  assign n972 = ~n803 & ~n971;
  assign n973 = ~n801 & n972;
  assign n974 = ~n796 & n973;
  assign n975 = ~n775 & n974;
  assign n976 = ~\in248  & \in348 ;
  assign n977 = ~\in255  & \in355 ;
  assign n978 = ~\in254  & \in354 ;
  assign n979 = ~n977 & ~n978;
  assign n980 = ~\in253  & \in353 ;
  assign n981 = ~\in252  & \in352 ;
  assign n982 = ~n980 & ~n981;
  assign n983 = n979 & n982;
  assign n984 = ~\in249  & \in349 ;
  assign n985 = ~\in251  & \in351 ;
  assign n986 = ~\in250  & \in350 ;
  assign n987 = ~n985 & ~n986;
  assign n988 = ~n984 & n987;
  assign n989 = n983 & n988;
  assign n990 = ~n976 & n989;
  assign n991 = ~n975 & n990;
  assign n992 = \in255  & ~\in355 ;
  assign n993 = \in251  & ~\in351 ;
  assign n994 = ~\in348  & ~n984;
  assign n995 = \in248  & n994;
  assign n996 = \in249  & ~\in349 ;
  assign n997 = ~n995 & ~n996;
  assign n998 = \in250  & ~\in350 ;
  assign n999 = n997 & ~n998;
  assign n1000 = n987 & ~n999;
  assign n1001 = ~n993 & ~n1000;
  assign n1002 = n983 & ~n1001;
  assign n1003 = \in252  & ~\in352 ;
  assign n1004 = ~n980 & n1003;
  assign n1005 = \in253  & ~\in353 ;
  assign n1006 = ~n1004 & ~n1005;
  assign n1007 = \in254  & ~\in354 ;
  assign n1008 = n1006 & ~n1007;
  assign n1009 = n979 & ~n1008;
  assign n1010 = ~n1002 & ~n1009;
  assign n1011 = ~n992 & n1010;
  assign n1012 = ~n991 & n1011;
  assign n1013 = ~\in256  & \in356 ;
  assign n1014 = ~n758 & ~n1013;
  assign n1015 = n753 & n1014;
  assign n1016 = n757 & n1015;
  assign n1017 = ~n1012 & n1016;
  assign n1018 = ~n774 & ~n1017;
  assign n1019 = ~n772 & n1018;
  assign n1020 = ~n767 & n1019;
  assign n1021 = ~n746 & n1020;
  assign n1022 = ~\in264  & \in364 ;
  assign n1023 = ~n1021 & ~n1022;
  assign n1024 = ~n745 & n1023;
  assign n1025 = n744 & n1024;
  assign n1026 = \in267  & ~\in367 ;
  assign n1027 = \in264  & ~\in364 ;
  assign n1028 = ~n745 & n1027;
  assign n1029 = \in265  & ~\in365 ;
  assign n1030 = ~n1028 & ~n1029;
  assign n1031 = \in266  & ~\in366 ;
  assign n1032 = n1030 & ~n1031;
  assign n1033 = n744 & ~n1032;
  assign n1034 = ~n1026 & ~n1033;
  assign n1035 = ~n1025 & n1034;
  assign n1036 = ~\in268  & \in368 ;
  assign n1037 = ~n734 & ~n1036;
  assign n1038 = n733 & n1037;
  assign n1039 = ~n1035 & n1038;
  assign n1040 = ~n741 & ~n1039;
  assign n1041 = ~n739 & n1040;
  assign n1042 = ~n730 & n1041;
  assign n1043 = ~\in275  & \in375 ;
  assign n1044 = ~\in274  & \in374 ;
  assign n1045 = ~n1043 & ~n1044;
  assign n1046 = ~\in273  & \in373 ;
  assign n1047 = ~\in272  & \in372 ;
  assign n1048 = ~n1046 & ~n1047;
  assign n1049 = n1045 & n1048;
  assign n1050 = ~n1042 & n1049;
  assign n1051 = \in275  & ~\in375 ;
  assign n1052 = \in272  & ~\in372 ;
  assign n1053 = ~n1046 & n1052;
  assign n1054 = \in273  & ~\in373 ;
  assign n1055 = ~n1053 & ~n1054;
  assign n1056 = \in274  & ~\in374 ;
  assign n1057 = n1055 & ~n1056;
  assign n1058 = n1045 & ~n1057;
  assign n1059 = ~n1051 & ~n1058;
  assign n1060 = ~n1050 & n1059;
  assign n1061 = ~\in276  & \in376 ;
  assign n1062 = ~n722 & ~n1061;
  assign n1063 = n721 & n1062;
  assign n1064 = ~n1060 & n1063;
  assign n1065 = ~n729 & ~n1064;
  assign n1066 = ~n727 & n1065;
  assign n1067 = ~n718 & n1066;
  assign n1068 = ~n717 & ~n1067;
  assign n1069 = n716 & n1068;
  assign n1070 = ~n713 & n1069;
  assign n1071 = \in283  & ~\in383 ;
  assign n1072 = ~\in380  & ~n717;
  assign n1073 = \in280  & n1072;
  assign n1074 = \in281  & ~\in381 ;
  assign n1075 = ~n1073 & ~n1074;
  assign n1076 = \in282  & ~\in382 ;
  assign n1077 = n1075 & ~n1076;
  assign n1078 = n716 & ~n1077;
  assign n1079 = ~n1071 & ~n1078;
  assign n1080 = ~n1070 & n1079;
  assign n1081 = ~\in284  & \in384 ;
  assign n1082 = ~n705 & ~n1081;
  assign n1083 = n704 & n1082;
  assign n1084 = ~n1080 & n1083;
  assign n1085 = ~n712 & ~n1084;
  assign n1086 = ~n710 & n1085;
  assign n1087 = ~n701 & n1086;
  assign n1088 = ~\in291  & \in391 ;
  assign n1089 = ~\in290  & \in390 ;
  assign n1090 = ~n1088 & ~n1089;
  assign n1091 = ~\in289  & \in389 ;
  assign n1092 = ~\in288  & \in388 ;
  assign n1093 = ~n1091 & ~n1092;
  assign n1094 = n1090 & n1093;
  assign n1095 = ~n1087 & n1094;
  assign n1096 = \in291  & ~\in391 ;
  assign n1097 = \in288  & ~\in388 ;
  assign n1098 = ~n1091 & n1097;
  assign n1099 = \in289  & ~\in389 ;
  assign n1100 = ~n1098 & ~n1099;
  assign n1101 = \in290  & ~\in390 ;
  assign n1102 = n1100 & ~n1101;
  assign n1103 = n1090 & ~n1102;
  assign n1104 = ~n1096 & ~n1103;
  assign n1105 = ~n1095 & n1104;
  assign n1106 = ~\in292  & \in392 ;
  assign n1107 = ~n693 & ~n1106;
  assign n1108 = n692 & n1107;
  assign n1109 = ~n1105 & n1108;
  assign n1110 = ~n700 & ~n1109;
  assign n1111 = ~n698 & n1110;
  assign n1112 = ~n689 & n1111;
  assign n1113 = ~n688 & ~n1112;
  assign n1114 = n687 & n1113;
  assign n1115 = ~n684 & n1114;
  assign n1116 = \in299  & ~\in399 ;
  assign n1117 = ~\in396  & ~n688;
  assign n1118 = \in296  & n1117;
  assign n1119 = \in297  & ~\in397 ;
  assign n1120 = ~n1118 & ~n1119;
  assign n1121 = \in298  & ~\in398 ;
  assign n1122 = n1120 & ~n1121;
  assign n1123 = n687 & ~n1122;
  assign n1124 = ~n1116 & ~n1123;
  assign n1125 = ~n1115 & n1124;
  assign n1126 = ~\in2100  & \in3100 ;
  assign n1127 = ~n676 & ~n1126;
  assign n1128 = n675 & n1127;
  assign n1129 = ~n1125 & n1128;
  assign n1130 = ~n683 & ~n1129;
  assign n1131 = ~n681 & n1130;
  assign n1132 = ~n672 & n1131;
  assign n1133 = ~\in2107  & \in3107 ;
  assign n1134 = ~\in2106  & \in3106 ;
  assign n1135 = ~n1133 & ~n1134;
  assign n1136 = ~\in2105  & \in3105 ;
  assign n1137 = ~\in2104  & \in3104 ;
  assign n1138 = ~n1136 & ~n1137;
  assign n1139 = n1135 & n1138;
  assign n1140 = ~n1132 & n1139;
  assign n1141 = \in2107  & ~\in3107 ;
  assign n1142 = \in2104  & ~\in3104 ;
  assign n1143 = ~n1136 & n1142;
  assign n1144 = \in2105  & ~\in3105 ;
  assign n1145 = ~n1143 & ~n1144;
  assign n1146 = \in2106  & ~\in3106 ;
  assign n1147 = n1145 & ~n1146;
  assign n1148 = n1135 & ~n1147;
  assign n1149 = ~n1141 & ~n1148;
  assign n1150 = ~n1140 & n1149;
  assign n1151 = ~\in2108  & \in3108 ;
  assign n1152 = ~n664 & ~n1151;
  assign n1153 = n663 & n1152;
  assign n1154 = ~n1150 & n1153;
  assign n1155 = ~n671 & ~n1154;
  assign n1156 = ~n669 & n1155;
  assign n1157 = ~n660 & n1156;
  assign n1158 = ~n659 & ~n1157;
  assign n1159 = n658 & n1158;
  assign n1160 = ~n655 & n1159;
  assign n1161 = \in2115  & ~\in3115 ;
  assign n1162 = ~\in3112  & ~n659;
  assign n1163 = \in2112  & n1162;
  assign n1164 = \in2113  & ~\in3113 ;
  assign n1165 = ~n1163 & ~n1164;
  assign n1166 = \in2114  & ~\in3114 ;
  assign n1167 = n1165 & ~n1166;
  assign n1168 = n658 & ~n1167;
  assign n1169 = ~n1161 & ~n1168;
  assign n1170 = ~n1160 & n1169;
  assign n1171 = ~\in2116  & \in3116 ;
  assign n1172 = ~n647 & ~n1171;
  assign n1173 = n646 & n1172;
  assign n1174 = ~n1170 & n1173;
  assign n1175 = ~n654 & ~n1174;
  assign n1176 = ~n652 & n1175;
  assign n1177 = ~n643 & n1176;
  assign n1178 = ~\in2123  & \in3123 ;
  assign n1179 = ~\in2122  & \in3122 ;
  assign n1180 = ~n1178 & ~n1179;
  assign n1181 = ~\in2121  & \in3121 ;
  assign n1182 = ~\in2120  & \in3120 ;
  assign n1183 = ~n1181 & ~n1182;
  assign n1184 = n1180 & n1183;
  assign n1185 = ~n1177 & n1184;
  assign n1186 = \in2123  & ~\in3123 ;
  assign n1187 = \in2120  & ~\in3120 ;
  assign n1188 = ~n1181 & n1187;
  assign n1189 = \in2121  & ~\in3121 ;
  assign n1190 = ~n1188 & ~n1189;
  assign n1191 = \in2122  & ~\in3122 ;
  assign n1192 = n1190 & ~n1191;
  assign n1193 = n1180 & ~n1192;
  assign n1194 = ~n1186 & ~n1193;
  assign n1195 = ~n1185 & n1194;
  assign n1196 = ~\in2124  & \in3124 ;
  assign n1197 = \in2127  & ~\in3127 ;
  assign n1198 = ~\in2126  & \in3126 ;
  assign n1199 = ~\in2125  & \in3125 ;
  assign n1200 = ~n1198 & ~n1199;
  assign n1201 = ~n1197 & n1200;
  assign n1202 = ~n1196 & n1201;
  assign n1203 = ~n1195 & n1202;
  assign n1204 = \in2124  & ~\in3124 ;
  assign n1205 = \in2125  & ~\in3125 ;
  assign n1206 = ~n1204 & ~n1205;
  assign n1207 = n1200 & ~n1206;
  assign n1208 = \in2126  & ~\in3126 ;
  assign n1209 = ~n1207 & ~n1208;
  assign n1210 = ~n1197 & ~n1209;
  assign n1211 = ~n1203 & ~n1210;
  assign n1212 = ~\in3127  & n1211;
  assign n1213 = \in2127  & ~n1212;
  assign n1214 = \in0119  & ~\in1119 ;
  assign n1215 = ~\in0119  & \in1119 ;
  assign n1216 = ~\in0118  & \in1118 ;
  assign n1217 = ~n1215 & ~n1216;
  assign n1218 = ~\in0117  & \in1117 ;
  assign n1219 = \in0116  & ~\in1116 ;
  assign n1220 = ~n1218 & n1219;
  assign n1221 = \in0117  & ~\in1117 ;
  assign n1222 = ~n1220 & ~n1221;
  assign n1223 = n1217 & ~n1222;
  assign n1224 = ~\in1118  & ~n1215;
  assign n1225 = \in0118  & n1224;
  assign n1226 = ~\in0112  & \in1112 ;
  assign n1227 = ~\in0115  & \in1115 ;
  assign n1228 = ~\in0114  & \in1114 ;
  assign n1229 = ~n1227 & ~n1228;
  assign n1230 = ~\in0113  & \in1113 ;
  assign n1231 = \in0111  & ~\in1111 ;
  assign n1232 = ~\in0111  & \in1111 ;
  assign n1233 = ~\in0110  & \in1110 ;
  assign n1234 = ~n1232 & ~n1233;
  assign n1235 = ~\in0109  & \in1109 ;
  assign n1236 = \in0108  & ~\in1108 ;
  assign n1237 = ~n1235 & n1236;
  assign n1238 = \in0109  & ~\in1109 ;
  assign n1239 = ~n1237 & ~n1238;
  assign n1240 = n1234 & ~n1239;
  assign n1241 = ~\in1110  & ~n1232;
  assign n1242 = \in0110  & n1241;
  assign n1243 = \in0103  & ~\in1103 ;
  assign n1244 = ~\in0103  & \in1103 ;
  assign n1245 = ~\in0102  & \in1102 ;
  assign n1246 = ~n1244 & ~n1245;
  assign n1247 = ~\in0101  & \in1101 ;
  assign n1248 = \in0100  & ~\in1100 ;
  assign n1249 = ~n1247 & n1248;
  assign n1250 = \in0101  & ~\in1101 ;
  assign n1251 = ~n1249 & ~n1250;
  assign n1252 = n1246 & ~n1251;
  assign n1253 = ~\in1102  & ~n1244;
  assign n1254 = \in0102  & n1253;
  assign n1255 = ~\in096  & \in196 ;
  assign n1256 = ~\in099  & \in199 ;
  assign n1257 = ~\in098  & \in198 ;
  assign n1258 = ~n1256 & ~n1257;
  assign n1259 = ~\in097  & \in197 ;
  assign n1260 = \in095  & ~\in195 ;
  assign n1261 = ~\in095  & \in195 ;
  assign n1262 = ~\in094  & \in194 ;
  assign n1263 = ~n1261 & ~n1262;
  assign n1264 = ~\in093  & \in193 ;
  assign n1265 = \in092  & ~\in192 ;
  assign n1266 = ~n1264 & n1265;
  assign n1267 = \in093  & ~\in193 ;
  assign n1268 = ~n1266 & ~n1267;
  assign n1269 = n1263 & ~n1268;
  assign n1270 = ~\in194  & ~n1261;
  assign n1271 = \in094  & n1270;
  assign n1272 = \in087  & ~\in187 ;
  assign n1273 = ~\in087  & \in187 ;
  assign n1274 = ~\in086  & \in186 ;
  assign n1275 = ~n1273 & ~n1274;
  assign n1276 = ~\in085  & \in185 ;
  assign n1277 = \in084  & ~\in184 ;
  assign n1278 = ~n1276 & n1277;
  assign n1279 = \in085  & ~\in185 ;
  assign n1280 = ~n1278 & ~n1279;
  assign n1281 = n1275 & ~n1280;
  assign n1282 = ~\in186  & ~n1273;
  assign n1283 = \in086  & n1282;
  assign n1284 = ~\in080  & \in180 ;
  assign n1285 = ~\in083  & \in183 ;
  assign n1286 = ~\in082  & \in182 ;
  assign n1287 = ~n1285 & ~n1286;
  assign n1288 = ~\in081  & \in181 ;
  assign n1289 = \in079  & ~\in179 ;
  assign n1290 = ~\in079  & \in179 ;
  assign n1291 = ~\in078  & \in178 ;
  assign n1292 = ~n1290 & ~n1291;
  assign n1293 = ~\in077  & \in177 ;
  assign n1294 = \in076  & ~\in176 ;
  assign n1295 = ~n1293 & n1294;
  assign n1296 = \in077  & ~\in177 ;
  assign n1297 = ~n1295 & ~n1296;
  assign n1298 = n1292 & ~n1297;
  assign n1299 = ~\in178  & ~n1290;
  assign n1300 = \in078  & n1299;
  assign n1301 = \in071  & ~\in171 ;
  assign n1302 = ~\in071  & \in171 ;
  assign n1303 = ~\in070  & \in170 ;
  assign n1304 = ~n1302 & ~n1303;
  assign n1305 = ~\in069  & \in169 ;
  assign n1306 = \in068  & ~\in168 ;
  assign n1307 = ~n1305 & n1306;
  assign n1308 = \in069  & ~\in169 ;
  assign n1309 = ~n1307 & ~n1308;
  assign n1310 = n1304 & ~n1309;
  assign n1311 = ~\in170  & ~n1302;
  assign n1312 = \in070  & n1311;
  assign n1313 = ~\in067  & \in167 ;
  assign n1314 = ~\in066  & \in166 ;
  assign n1315 = ~n1313 & ~n1314;
  assign n1316 = ~\in065  & \in165 ;
  assign n1317 = \in063  & ~\in163 ;
  assign n1318 = ~\in063  & \in163 ;
  assign n1319 = ~\in062  & \in162 ;
  assign n1320 = ~n1318 & ~n1319;
  assign n1321 = ~\in060  & \in160 ;
  assign n1322 = ~\in061  & \in161 ;
  assign n1323 = ~n1321 & ~n1322;
  assign n1324 = n1320 & n1323;
  assign n1325 = \in059  & ~\in159 ;
  assign n1326 = ~\in059  & \in159 ;
  assign n1327 = ~\in058  & \in158 ;
  assign n1328 = ~n1326 & ~n1327;
  assign n1329 = ~\in057  & \in157 ;
  assign n1330 = \in056  & ~\in156 ;
  assign n1331 = ~n1329 & n1330;
  assign n1332 = \in057  & ~\in157 ;
  assign n1333 = ~n1331 & ~n1332;
  assign n1334 = \in058  & ~\in158 ;
  assign n1335 = n1333 & ~n1334;
  assign n1336 = n1328 & ~n1335;
  assign n1337 = ~n1325 & ~n1336;
  assign n1338 = n1324 & ~n1337;
  assign n1339 = \in060  & ~\in160 ;
  assign n1340 = ~n1322 & n1339;
  assign n1341 = \in061  & ~\in161 ;
  assign n1342 = ~n1340 & ~n1341;
  assign n1343 = n1320 & ~n1342;
  assign n1344 = ~\in162  & ~n1318;
  assign n1345 = \in062  & n1344;
  assign n1346 = \in047  & ~\in147 ;
  assign n1347 = ~\in047  & \in147 ;
  assign n1348 = ~\in046  & \in146 ;
  assign n1349 = ~n1347 & ~n1348;
  assign n1350 = ~\in044  & \in144 ;
  assign n1351 = ~\in045  & \in145 ;
  assign n1352 = ~n1350 & ~n1351;
  assign n1353 = n1349 & n1352;
  assign n1354 = \in043  & ~\in143 ;
  assign n1355 = ~\in043  & \in143 ;
  assign n1356 = ~\in042  & \in142 ;
  assign n1357 = ~n1355 & ~n1356;
  assign n1358 = ~\in041  & \in141 ;
  assign n1359 = \in040  & ~\in140 ;
  assign n1360 = ~n1358 & n1359;
  assign n1361 = \in041  & ~\in141 ;
  assign n1362 = ~n1360 & ~n1361;
  assign n1363 = \in042  & ~\in142 ;
  assign n1364 = n1362 & ~n1363;
  assign n1365 = n1357 & ~n1364;
  assign n1366 = ~n1354 & ~n1365;
  assign n1367 = n1353 & ~n1366;
  assign n1368 = \in044  & ~\in144 ;
  assign n1369 = ~n1351 & n1368;
  assign n1370 = \in045  & ~\in145 ;
  assign n1371 = ~n1369 & ~n1370;
  assign n1372 = n1349 & ~n1371;
  assign n1373 = ~\in146  & ~n1347;
  assign n1374 = \in046  & n1373;
  assign n1375 = ~\in032  & \in132 ;
  assign n1376 = ~\in031  & \in131 ;
  assign n1377 = ~\in030  & \in130 ;
  assign n1378 = ~\in029  & \in129 ;
  assign n1379 = ~\in028  & \in128 ;
  assign n1380 = ~\in027  & \in127 ;
  assign n1381 = ~\in026  & \in126 ;
  assign n1382 = ~\in023  & \in123 ;
  assign n1383 = ~\in022  & \in122 ;
  assign n1384 = ~\in021  & \in121 ;
  assign n1385 = ~\in020  & \in120 ;
  assign n1386 = ~\in019  & \in119 ;
  assign n1387 = ~\in018  & \in118 ;
  assign n1388 = ~\in015  & \in115 ;
  assign n1389 = ~\in014  & \in114 ;
  assign n1390 = ~\in013  & \in113 ;
  assign n1391 = ~\in012  & \in112 ;
  assign n1392 = ~\in011  & \in111 ;
  assign n1393 = ~\in010  & \in110 ;
  assign n1394 = ~\in07  & \in17 ;
  assign n1395 = ~\in06  & \in16 ;
  assign n1396 = ~\in03  & \in13 ;
  assign n1397 = \in00  & ~\in10 ;
  assign n1398 = \in01  & ~\in11 ;
  assign n1399 = ~n1397 & ~n1398;
  assign n1400 = ~\in02  & \in12 ;
  assign n1401 = ~\in01  & \in11 ;
  assign n1402 = ~n1400 & ~n1401;
  assign n1403 = ~n1399 & n1402;
  assign n1404 = \in02  & ~\in12 ;
  assign n1405 = ~n1403 & ~n1404;
  assign n1406 = ~n1396 & ~n1405;
  assign n1407 = \in03  & ~\in13 ;
  assign n1408 = ~n1406 & ~n1407;
  assign n1409 = ~\in04  & n1408;
  assign n1410 = ~\in14  & ~n1409;
  assign n1411 = \in04  & ~n1408;
  assign n1412 = ~n1410 & ~n1411;
  assign n1413 = ~\in05  & n1412;
  assign n1414 = ~\in15  & ~n1413;
  assign n1415 = \in05  & ~n1412;
  assign n1416 = ~n1414 & ~n1415;
  assign n1417 = ~n1395 & ~n1416;
  assign n1418 = \in06  & ~\in16 ;
  assign n1419 = ~n1417 & ~n1418;
  assign n1420 = ~n1394 & ~n1419;
  assign n1421 = \in07  & ~\in17 ;
  assign n1422 = ~n1420 & ~n1421;
  assign n1423 = ~\in08  & n1422;
  assign n1424 = ~\in18  & ~n1423;
  assign n1425 = \in08  & ~n1422;
  assign n1426 = ~n1424 & ~n1425;
  assign n1427 = ~\in09  & n1426;
  assign n1428 = ~\in19  & ~n1427;
  assign n1429 = \in09  & ~n1426;
  assign n1430 = ~n1428 & ~n1429;
  assign n1431 = ~n1393 & ~n1430;
  assign n1432 = \in010  & ~\in110 ;
  assign n1433 = ~n1431 & ~n1432;
  assign n1434 = ~n1392 & ~n1433;
  assign n1435 = \in011  & ~\in111 ;
  assign n1436 = ~n1434 & ~n1435;
  assign n1437 = ~n1391 & ~n1436;
  assign n1438 = \in012  & ~\in112 ;
  assign n1439 = ~n1437 & ~n1438;
  assign n1440 = ~n1390 & ~n1439;
  assign n1441 = \in013  & ~\in113 ;
  assign n1442 = ~n1440 & ~n1441;
  assign n1443 = ~n1389 & ~n1442;
  assign n1444 = \in014  & ~\in114 ;
  assign n1445 = ~n1443 & ~n1444;
  assign n1446 = ~n1388 & ~n1445;
  assign n1447 = \in015  & ~\in115 ;
  assign n1448 = ~n1446 & ~n1447;
  assign n1449 = ~\in016  & n1448;
  assign n1450 = ~\in116  & ~n1449;
  assign n1451 = \in016  & ~n1448;
  assign n1452 = ~n1450 & ~n1451;
  assign n1453 = ~\in017  & n1452;
  assign n1454 = ~\in117  & ~n1453;
  assign n1455 = \in017  & ~n1452;
  assign n1456 = ~n1454 & ~n1455;
  assign n1457 = ~n1387 & ~n1456;
  assign n1458 = \in018  & ~\in118 ;
  assign n1459 = ~n1457 & ~n1458;
  assign n1460 = ~n1386 & ~n1459;
  assign n1461 = \in019  & ~\in119 ;
  assign n1462 = ~n1460 & ~n1461;
  assign n1463 = ~n1385 & ~n1462;
  assign n1464 = \in020  & ~\in120 ;
  assign n1465 = ~n1463 & ~n1464;
  assign n1466 = ~n1384 & ~n1465;
  assign n1467 = \in021  & ~\in121 ;
  assign n1468 = ~n1466 & ~n1467;
  assign n1469 = ~n1383 & ~n1468;
  assign n1470 = \in022  & ~\in122 ;
  assign n1471 = ~n1469 & ~n1470;
  assign n1472 = ~n1382 & ~n1471;
  assign n1473 = \in023  & ~\in123 ;
  assign n1474 = ~n1472 & ~n1473;
  assign n1475 = ~\in024  & n1474;
  assign n1476 = ~\in124  & ~n1475;
  assign n1477 = \in024  & ~n1474;
  assign n1478 = ~n1476 & ~n1477;
  assign n1479 = ~\in025  & n1478;
  assign n1480 = ~\in125  & ~n1479;
  assign n1481 = \in025  & ~n1478;
  assign n1482 = ~n1480 & ~n1481;
  assign n1483 = ~n1381 & ~n1482;
  assign n1484 = \in026  & ~\in126 ;
  assign n1485 = ~n1483 & ~n1484;
  assign n1486 = ~n1380 & ~n1485;
  assign n1487 = \in027  & ~\in127 ;
  assign n1488 = ~n1486 & ~n1487;
  assign n1489 = ~n1379 & ~n1488;
  assign n1490 = \in028  & ~\in128 ;
  assign n1491 = ~n1489 & ~n1490;
  assign n1492 = ~n1378 & ~n1491;
  assign n1493 = \in029  & ~\in129 ;
  assign n1494 = ~n1492 & ~n1493;
  assign n1495 = ~n1377 & ~n1494;
  assign n1496 = \in030  & ~\in130 ;
  assign n1497 = ~n1495 & ~n1496;
  assign n1498 = ~n1376 & ~n1497;
  assign n1499 = \in031  & ~\in131 ;
  assign n1500 = ~n1498 & ~n1499;
  assign n1501 = ~\in039  & \in139 ;
  assign n1502 = ~\in038  & \in138 ;
  assign n1503 = ~n1501 & ~n1502;
  assign n1504 = ~\in036  & \in136 ;
  assign n1505 = ~\in037  & \in137 ;
  assign n1506 = ~n1504 & ~n1505;
  assign n1507 = n1503 & n1506;
  assign n1508 = ~\in033  & \in133 ;
  assign n1509 = ~\in035  & \in135 ;
  assign n1510 = ~\in034  & \in134 ;
  assign n1511 = ~n1509 & ~n1510;
  assign n1512 = ~n1508 & n1511;
  assign n1513 = n1507 & n1512;
  assign n1514 = ~n1500 & n1513;
  assign n1515 = ~n1375 & n1514;
  assign n1516 = \in039  & ~\in139 ;
  assign n1517 = \in036  & ~\in136 ;
  assign n1518 = ~n1505 & n1517;
  assign n1519 = \in037  & ~\in137 ;
  assign n1520 = ~n1518 & ~n1519;
  assign n1521 = n1503 & ~n1520;
  assign n1522 = ~\in138  & ~n1501;
  assign n1523 = \in038  & n1522;
  assign n1524 = \in035  & ~\in135 ;
  assign n1525 = ~\in132  & ~n1508;
  assign n1526 = \in032  & n1525;
  assign n1527 = \in033  & ~\in133 ;
  assign n1528 = ~n1526 & ~n1527;
  assign n1529 = \in034  & ~\in134 ;
  assign n1530 = n1528 & ~n1529;
  assign n1531 = n1511 & ~n1530;
  assign n1532 = ~n1524 & ~n1531;
  assign n1533 = n1507 & ~n1532;
  assign n1534 = ~n1523 & ~n1533;
  assign n1535 = ~n1521 & n1534;
  assign n1536 = ~n1516 & n1535;
  assign n1537 = ~n1515 & n1536;
  assign n1538 = ~\in040  & \in140 ;
  assign n1539 = ~n1358 & ~n1538;
  assign n1540 = n1357 & n1539;
  assign n1541 = n1353 & n1540;
  assign n1542 = ~n1537 & n1541;
  assign n1543 = ~n1374 & ~n1542;
  assign n1544 = ~n1372 & n1543;
  assign n1545 = ~n1367 & n1544;
  assign n1546 = ~n1346 & n1545;
  assign n1547 = ~\in048  & \in148 ;
  assign n1548 = ~\in055  & \in155 ;
  assign n1549 = ~\in054  & \in154 ;
  assign n1550 = ~n1548 & ~n1549;
  assign n1551 = ~\in053  & \in153 ;
  assign n1552 = ~\in052  & \in152 ;
  assign n1553 = ~n1551 & ~n1552;
  assign n1554 = n1550 & n1553;
  assign n1555 = ~\in049  & \in149 ;
  assign n1556 = ~\in051  & \in151 ;
  assign n1557 = ~\in050  & \in150 ;
  assign n1558 = ~n1556 & ~n1557;
  assign n1559 = ~n1555 & n1558;
  assign n1560 = n1554 & n1559;
  assign n1561 = ~n1547 & n1560;
  assign n1562 = ~n1546 & n1561;
  assign n1563 = \in055  & ~\in155 ;
  assign n1564 = \in051  & ~\in151 ;
  assign n1565 = ~\in148  & ~n1555;
  assign n1566 = \in048  & n1565;
  assign n1567 = \in049  & ~\in149 ;
  assign n1568 = ~n1566 & ~n1567;
  assign n1569 = \in050  & ~\in150 ;
  assign n1570 = n1568 & ~n1569;
  assign n1571 = n1558 & ~n1570;
  assign n1572 = ~n1564 & ~n1571;
  assign n1573 = n1554 & ~n1572;
  assign n1574 = \in052  & ~\in152 ;
  assign n1575 = ~n1551 & n1574;
  assign n1576 = \in053  & ~\in153 ;
  assign n1577 = ~n1575 & ~n1576;
  assign n1578 = \in054  & ~\in154 ;
  assign n1579 = n1577 & ~n1578;
  assign n1580 = n1550 & ~n1579;
  assign n1581 = ~n1573 & ~n1580;
  assign n1582 = ~n1563 & n1581;
  assign n1583 = ~n1562 & n1582;
  assign n1584 = ~\in056  & \in156 ;
  assign n1585 = ~n1329 & ~n1584;
  assign n1586 = n1324 & n1585;
  assign n1587 = n1328 & n1586;
  assign n1588 = ~n1583 & n1587;
  assign n1589 = ~n1345 & ~n1588;
  assign n1590 = ~n1343 & n1589;
  assign n1591 = ~n1338 & n1590;
  assign n1592 = ~n1317 & n1591;
  assign n1593 = ~\in064  & \in164 ;
  assign n1594 = ~n1592 & ~n1593;
  assign n1595 = ~n1316 & n1594;
  assign n1596 = n1315 & n1595;
  assign n1597 = \in067  & ~\in167 ;
  assign n1598 = \in064  & ~\in164 ;
  assign n1599 = ~n1316 & n1598;
  assign n1600 = \in065  & ~\in165 ;
  assign n1601 = ~n1599 & ~n1600;
  assign n1602 = \in066  & ~\in166 ;
  assign n1603 = n1601 & ~n1602;
  assign n1604 = n1315 & ~n1603;
  assign n1605 = ~n1597 & ~n1604;
  assign n1606 = ~n1596 & n1605;
  assign n1607 = ~\in068  & \in168 ;
  assign n1608 = ~n1305 & ~n1607;
  assign n1609 = n1304 & n1608;
  assign n1610 = ~n1606 & n1609;
  assign n1611 = ~n1312 & ~n1610;
  assign n1612 = ~n1310 & n1611;
  assign n1613 = ~n1301 & n1612;
  assign n1614 = ~\in075  & \in175 ;
  assign n1615 = ~\in074  & \in174 ;
  assign n1616 = ~n1614 & ~n1615;
  assign n1617 = ~\in073  & \in173 ;
  assign n1618 = ~\in072  & \in172 ;
  assign n1619 = ~n1617 & ~n1618;
  assign n1620 = n1616 & n1619;
  assign n1621 = ~n1613 & n1620;
  assign n1622 = \in075  & ~\in175 ;
  assign n1623 = \in072  & ~\in172 ;
  assign n1624 = ~n1617 & n1623;
  assign n1625 = \in073  & ~\in173 ;
  assign n1626 = ~n1624 & ~n1625;
  assign n1627 = \in074  & ~\in174 ;
  assign n1628 = n1626 & ~n1627;
  assign n1629 = n1616 & ~n1628;
  assign n1630 = ~n1622 & ~n1629;
  assign n1631 = ~n1621 & n1630;
  assign n1632 = ~\in076  & \in176 ;
  assign n1633 = ~n1293 & ~n1632;
  assign n1634 = n1292 & n1633;
  assign n1635 = ~n1631 & n1634;
  assign n1636 = ~n1300 & ~n1635;
  assign n1637 = ~n1298 & n1636;
  assign n1638 = ~n1289 & n1637;
  assign n1639 = ~n1288 & ~n1638;
  assign n1640 = n1287 & n1639;
  assign n1641 = ~n1284 & n1640;
  assign n1642 = \in083  & ~\in183 ;
  assign n1643 = ~\in180  & ~n1288;
  assign n1644 = \in080  & n1643;
  assign n1645 = \in081  & ~\in181 ;
  assign n1646 = ~n1644 & ~n1645;
  assign n1647 = \in082  & ~\in182 ;
  assign n1648 = n1646 & ~n1647;
  assign n1649 = n1287 & ~n1648;
  assign n1650 = ~n1642 & ~n1649;
  assign n1651 = ~n1641 & n1650;
  assign n1652 = ~\in084  & \in184 ;
  assign n1653 = ~n1276 & ~n1652;
  assign n1654 = n1275 & n1653;
  assign n1655 = ~n1651 & n1654;
  assign n1656 = ~n1283 & ~n1655;
  assign n1657 = ~n1281 & n1656;
  assign n1658 = ~n1272 & n1657;
  assign n1659 = ~\in091  & \in191 ;
  assign n1660 = ~\in090  & \in190 ;
  assign n1661 = ~n1659 & ~n1660;
  assign n1662 = ~\in089  & \in189 ;
  assign n1663 = ~\in088  & \in188 ;
  assign n1664 = ~n1662 & ~n1663;
  assign n1665 = n1661 & n1664;
  assign n1666 = ~n1658 & n1665;
  assign n1667 = \in091  & ~\in191 ;
  assign n1668 = \in088  & ~\in188 ;
  assign n1669 = ~n1662 & n1668;
  assign n1670 = \in089  & ~\in189 ;
  assign n1671 = ~n1669 & ~n1670;
  assign n1672 = \in090  & ~\in190 ;
  assign n1673 = n1671 & ~n1672;
  assign n1674 = n1661 & ~n1673;
  assign n1675 = ~n1667 & ~n1674;
  assign n1676 = ~n1666 & n1675;
  assign n1677 = ~\in092  & \in192 ;
  assign n1678 = ~n1264 & ~n1677;
  assign n1679 = n1263 & n1678;
  assign n1680 = ~n1676 & n1679;
  assign n1681 = ~n1271 & ~n1680;
  assign n1682 = ~n1269 & n1681;
  assign n1683 = ~n1260 & n1682;
  assign n1684 = ~n1259 & ~n1683;
  assign n1685 = n1258 & n1684;
  assign n1686 = ~n1255 & n1685;
  assign n1687 = \in099  & ~\in199 ;
  assign n1688 = ~\in196  & ~n1259;
  assign n1689 = \in096  & n1688;
  assign n1690 = \in097  & ~\in197 ;
  assign n1691 = ~n1689 & ~n1690;
  assign n1692 = \in098  & ~\in198 ;
  assign n1693 = n1691 & ~n1692;
  assign n1694 = n1258 & ~n1693;
  assign n1695 = ~n1687 & ~n1694;
  assign n1696 = ~n1686 & n1695;
  assign n1697 = ~\in0100  & \in1100 ;
  assign n1698 = ~n1247 & ~n1697;
  assign n1699 = n1246 & n1698;
  assign n1700 = ~n1696 & n1699;
  assign n1701 = ~n1254 & ~n1700;
  assign n1702 = ~n1252 & n1701;
  assign n1703 = ~n1243 & n1702;
  assign n1704 = ~\in0107  & \in1107 ;
  assign n1705 = ~\in0106  & \in1106 ;
  assign n1706 = ~n1704 & ~n1705;
  assign n1707 = ~\in0105  & \in1105 ;
  assign n1708 = ~\in0104  & \in1104 ;
  assign n1709 = ~n1707 & ~n1708;
  assign n1710 = n1706 & n1709;
  assign n1711 = ~n1703 & n1710;
  assign n1712 = \in0107  & ~\in1107 ;
  assign n1713 = \in0104  & ~\in1104 ;
  assign n1714 = ~n1707 & n1713;
  assign n1715 = \in0105  & ~\in1105 ;
  assign n1716 = ~n1714 & ~n1715;
  assign n1717 = \in0106  & ~\in1106 ;
  assign n1718 = n1716 & ~n1717;
  assign n1719 = n1706 & ~n1718;
  assign n1720 = ~n1712 & ~n1719;
  assign n1721 = ~n1711 & n1720;
  assign n1722 = ~\in0108  & \in1108 ;
  assign n1723 = ~n1235 & ~n1722;
  assign n1724 = n1234 & n1723;
  assign n1725 = ~n1721 & n1724;
  assign n1726 = ~n1242 & ~n1725;
  assign n1727 = ~n1240 & n1726;
  assign n1728 = ~n1231 & n1727;
  assign n1729 = ~n1230 & ~n1728;
  assign n1730 = n1229 & n1729;
  assign n1731 = ~n1226 & n1730;
  assign n1732 = \in0115  & ~\in1115 ;
  assign n1733 = ~\in1112  & ~n1230;
  assign n1734 = \in0112  & n1733;
  assign n1735 = \in0113  & ~\in1113 ;
  assign n1736 = ~n1734 & ~n1735;
  assign n1737 = \in0114  & ~\in1114 ;
  assign n1738 = n1736 & ~n1737;
  assign n1739 = n1229 & ~n1738;
  assign n1740 = ~n1732 & ~n1739;
  assign n1741 = ~n1731 & n1740;
  assign n1742 = ~\in0116  & \in1116 ;
  assign n1743 = ~n1218 & ~n1742;
  assign n1744 = n1217 & n1743;
  assign n1745 = ~n1741 & n1744;
  assign n1746 = ~n1225 & ~n1745;
  assign n1747 = ~n1223 & n1746;
  assign n1748 = ~n1214 & n1747;
  assign n1749 = ~\in0123  & \in1123 ;
  assign n1750 = ~\in0122  & \in1122 ;
  assign n1751 = ~n1749 & ~n1750;
  assign n1752 = ~\in0121  & \in1121 ;
  assign n1753 = ~\in0120  & \in1120 ;
  assign n1754 = ~n1752 & ~n1753;
  assign n1755 = n1751 & n1754;
  assign n1756 = ~n1748 & n1755;
  assign n1757 = \in0123  & ~\in1123 ;
  assign n1758 = \in0120  & ~\in1120 ;
  assign n1759 = ~n1752 & n1758;
  assign n1760 = \in0121  & ~\in1121 ;
  assign n1761 = ~n1759 & ~n1760;
  assign n1762 = \in0122  & ~\in1122 ;
  assign n1763 = n1761 & ~n1762;
  assign n1764 = n1751 & ~n1763;
  assign n1765 = ~n1757 & ~n1764;
  assign n1766 = ~n1756 & n1765;
  assign n1767 = ~\in0124  & \in1124 ;
  assign n1768 = \in0127  & ~\in1127 ;
  assign n1769 = ~\in0126  & \in1126 ;
  assign n1770 = ~\in0125  & \in1125 ;
  assign n1771 = ~n1769 & ~n1770;
  assign n1772 = ~n1768 & n1771;
  assign n1773 = ~n1767 & n1772;
  assign n1774 = ~n1766 & n1773;
  assign n1775 = \in0124  & ~\in1124 ;
  assign n1776 = \in0125  & ~\in1125 ;
  assign n1777 = ~n1775 & ~n1776;
  assign n1778 = n1771 & ~n1777;
  assign n1779 = \in0126  & ~\in1126 ;
  assign n1780 = ~n1778 & ~n1779;
  assign n1781 = ~n1768 & ~n1780;
  assign n1782 = ~n1774 & ~n1781;
  assign n1783 = ~\in1127  & n1782;
  assign n1784 = \in0127  & ~n1783;
  assign n1785 = n1213 & ~n1784;
  assign n1786 = ~\in0127  & \in1127 ;
  assign n1787 = n1782 & ~n1786;
  assign n1788 = \in1119  & n1787;
  assign n1789 = \in0119  & ~n1787;
  assign n1790 = ~n1788 & ~n1789;
  assign n1791 = ~\in2127  & \in3127 ;
  assign n1792 = n1211 & ~n1791;
  assign n1793 = \in3119  & n1792;
  assign n1794 = \in2119  & ~n1792;
  assign n1795 = ~n1793 & ~n1794;
  assign n1796 = ~n1790 & n1795;
  assign n1797 = n1790 & ~n1795;
  assign n1798 = \in3118  & n1792;
  assign n1799 = \in2118  & ~n1792;
  assign n1800 = ~n1798 & ~n1799;
  assign n1801 = \in1118  & n1787;
  assign n1802 = \in0118  & ~n1787;
  assign n1803 = ~n1801 & ~n1802;
  assign n1804 = ~n1800 & n1803;
  assign n1805 = ~n1797 & ~n1804;
  assign n1806 = \in1116  & n1787;
  assign n1807 = \in0116  & ~n1787;
  assign n1808 = ~n1806 & ~n1807;
  assign n1809 = \in1117  & n1787;
  assign n1810 = \in0117  & ~n1787;
  assign n1811 = ~n1809 & ~n1810;
  assign n1812 = \in3117  & n1792;
  assign n1813 = \in2117  & ~n1792;
  assign n1814 = ~n1812 & ~n1813;
  assign n1815 = n1811 & ~n1814;
  assign n1816 = \in3116  & n1792;
  assign n1817 = \in2116  & ~n1792;
  assign n1818 = ~n1816 & ~n1817;
  assign n1819 = ~n1815 & n1818;
  assign n1820 = ~n1808 & n1819;
  assign n1821 = ~n1811 & n1814;
  assign n1822 = ~n1820 & ~n1821;
  assign n1823 = n1805 & ~n1822;
  assign n1824 = n1800 & ~n1803;
  assign n1825 = ~n1797 & n1824;
  assign n1826 = \in3112  & n1792;
  assign n1827 = \in2112  & ~n1792;
  assign n1828 = ~n1826 & ~n1827;
  assign n1829 = \in1112  & n1787;
  assign n1830 = \in0112  & ~n1787;
  assign n1831 = ~n1829 & ~n1830;
  assign n1832 = ~n1828 & n1831;
  assign n1833 = \in1115  & n1787;
  assign n1834 = \in0115  & ~n1787;
  assign n1835 = ~n1833 & ~n1834;
  assign n1836 = \in3115  & n1792;
  assign n1837 = \in2115  & ~n1792;
  assign n1838 = ~n1836 & ~n1837;
  assign n1839 = n1835 & ~n1838;
  assign n1840 = \in3114  & n1792;
  assign n1841 = \in2114  & ~n1792;
  assign n1842 = ~n1840 & ~n1841;
  assign n1843 = \in1114  & n1787;
  assign n1844 = \in0114  & ~n1787;
  assign n1845 = ~n1843 & ~n1844;
  assign n1846 = ~n1842 & n1845;
  assign n1847 = ~n1839 & ~n1846;
  assign n1848 = \in1113  & n1787;
  assign n1849 = \in0113  & ~n1787;
  assign n1850 = ~n1848 & ~n1849;
  assign n1851 = \in3113  & n1792;
  assign n1852 = \in2113  & ~n1792;
  assign n1853 = ~n1851 & ~n1852;
  assign n1854 = n1850 & ~n1853;
  assign n1855 = \in1111  & n1787;
  assign n1856 = \in0111  & ~n1787;
  assign n1857 = ~n1855 & ~n1856;
  assign n1858 = \in3111  & n1792;
  assign n1859 = \in2111  & ~n1792;
  assign n1860 = ~n1858 & ~n1859;
  assign n1861 = ~n1857 & n1860;
  assign n1862 = n1857 & ~n1860;
  assign n1863 = \in3110  & n1792;
  assign n1864 = \in2110  & ~n1792;
  assign n1865 = ~n1863 & ~n1864;
  assign n1866 = \in1110  & n1787;
  assign n1867 = \in0110  & ~n1787;
  assign n1868 = ~n1866 & ~n1867;
  assign n1869 = ~n1865 & n1868;
  assign n1870 = ~n1862 & ~n1869;
  assign n1871 = \in1109  & n1787;
  assign n1872 = \in0109  & ~n1787;
  assign n1873 = ~n1871 & ~n1872;
  assign n1874 = \in3109  & n1792;
  assign n1875 = \in2109  & ~n1792;
  assign n1876 = ~n1874 & ~n1875;
  assign n1877 = n1873 & ~n1876;
  assign n1878 = \in1108  & n1787;
  assign n1879 = \in0108  & ~n1787;
  assign n1880 = ~n1878 & ~n1879;
  assign n1881 = \in3108  & n1792;
  assign n1882 = \in2108  & ~n1792;
  assign n1883 = ~n1881 & ~n1882;
  assign n1884 = ~n1880 & n1883;
  assign n1885 = ~n1877 & n1884;
  assign n1886 = ~n1873 & n1876;
  assign n1887 = ~n1885 & ~n1886;
  assign n1888 = n1870 & ~n1887;
  assign n1889 = n1865 & ~n1868;
  assign n1890 = ~n1862 & n1889;
  assign n1891 = \in1103  & n1787;
  assign n1892 = \in0103  & ~n1787;
  assign n1893 = ~n1891 & ~n1892;
  assign n1894 = \in3103  & n1792;
  assign n1895 = \in2103  & ~n1792;
  assign n1896 = ~n1894 & ~n1895;
  assign n1897 = ~n1893 & n1896;
  assign n1898 = n1893 & ~n1896;
  assign n1899 = \in3102  & n1792;
  assign n1900 = \in2102  & ~n1792;
  assign n1901 = ~n1899 & ~n1900;
  assign n1902 = \in1102  & n1787;
  assign n1903 = \in0102  & ~n1787;
  assign n1904 = ~n1902 & ~n1903;
  assign n1905 = ~n1901 & n1904;
  assign n1906 = ~n1898 & ~n1905;
  assign n1907 = \in1101  & n1787;
  assign n1908 = \in0101  & ~n1787;
  assign n1909 = ~n1907 & ~n1908;
  assign n1910 = \in3101  & n1792;
  assign n1911 = \in2101  & ~n1792;
  assign n1912 = ~n1910 & ~n1911;
  assign n1913 = n1909 & ~n1912;
  assign n1914 = \in1100  & n1787;
  assign n1915 = \in0100  & ~n1787;
  assign n1916 = ~n1914 & ~n1915;
  assign n1917 = \in3100  & n1792;
  assign n1918 = \in2100  & ~n1792;
  assign n1919 = ~n1917 & ~n1918;
  assign n1920 = ~n1916 & n1919;
  assign n1921 = ~n1913 & n1920;
  assign n1922 = ~n1909 & n1912;
  assign n1923 = ~n1921 & ~n1922;
  assign n1924 = n1906 & ~n1923;
  assign n1925 = n1901 & ~n1904;
  assign n1926 = ~n1898 & n1925;
  assign n1927 = \in396  & n1792;
  assign n1928 = \in296  & ~n1792;
  assign n1929 = ~n1927 & ~n1928;
  assign n1930 = \in196  & n1787;
  assign n1931 = \in096  & ~n1787;
  assign n1932 = ~n1930 & ~n1931;
  assign n1933 = ~n1929 & n1932;
  assign n1934 = \in199  & n1787;
  assign n1935 = \in099  & ~n1787;
  assign n1936 = ~n1934 & ~n1935;
  assign n1937 = \in399  & n1792;
  assign n1938 = \in299  & ~n1792;
  assign n1939 = ~n1937 & ~n1938;
  assign n1940 = n1936 & ~n1939;
  assign n1941 = \in398  & n1792;
  assign n1942 = \in298  & ~n1792;
  assign n1943 = ~n1941 & ~n1942;
  assign n1944 = \in198  & n1787;
  assign n1945 = \in098  & ~n1787;
  assign n1946 = ~n1944 & ~n1945;
  assign n1947 = ~n1943 & n1946;
  assign n1948 = ~n1940 & ~n1947;
  assign n1949 = \in197  & n1787;
  assign n1950 = \in097  & ~n1787;
  assign n1951 = ~n1949 & ~n1950;
  assign n1952 = \in397  & n1792;
  assign n1953 = \in297  & ~n1792;
  assign n1954 = ~n1952 & ~n1953;
  assign n1955 = n1951 & ~n1954;
  assign n1956 = \in195  & n1787;
  assign n1957 = \in095  & ~n1787;
  assign n1958 = ~n1956 & ~n1957;
  assign n1959 = \in395  & n1792;
  assign n1960 = \in295  & ~n1792;
  assign n1961 = ~n1959 & ~n1960;
  assign n1962 = ~n1958 & n1961;
  assign n1963 = n1958 & ~n1961;
  assign n1964 = \in394  & n1792;
  assign n1965 = \in294  & ~n1792;
  assign n1966 = ~n1964 & ~n1965;
  assign n1967 = \in194  & n1787;
  assign n1968 = \in094  & ~n1787;
  assign n1969 = ~n1967 & ~n1968;
  assign n1970 = ~n1966 & n1969;
  assign n1971 = ~n1963 & ~n1970;
  assign n1972 = \in193  & n1787;
  assign n1973 = \in093  & ~n1787;
  assign n1974 = ~n1972 & ~n1973;
  assign n1975 = \in393  & n1792;
  assign n1976 = \in293  & ~n1792;
  assign n1977 = ~n1975 & ~n1976;
  assign n1978 = n1974 & ~n1977;
  assign n1979 = \in192  & n1787;
  assign n1980 = \in092  & ~n1787;
  assign n1981 = ~n1979 & ~n1980;
  assign n1982 = \in392  & n1792;
  assign n1983 = \in292  & ~n1792;
  assign n1984 = ~n1982 & ~n1983;
  assign n1985 = ~n1981 & n1984;
  assign n1986 = ~n1978 & n1985;
  assign n1987 = ~n1974 & n1977;
  assign n1988 = ~n1986 & ~n1987;
  assign n1989 = n1971 & ~n1988;
  assign n1990 = n1966 & ~n1969;
  assign n1991 = ~n1963 & n1990;
  assign n1992 = \in187  & n1787;
  assign n1993 = \in087  & ~n1787;
  assign n1994 = ~n1992 & ~n1993;
  assign n1995 = \in387  & n1792;
  assign n1996 = \in287  & ~n1792;
  assign n1997 = ~n1995 & ~n1996;
  assign n1998 = ~n1994 & n1997;
  assign n1999 = n1994 & ~n1997;
  assign n2000 = \in386  & n1792;
  assign n2001 = \in286  & ~n1792;
  assign n2002 = ~n2000 & ~n2001;
  assign n2003 = \in186  & n1787;
  assign n2004 = \in086  & ~n1787;
  assign n2005 = ~n2003 & ~n2004;
  assign n2006 = ~n2002 & n2005;
  assign n2007 = ~n1999 & ~n2006;
  assign n2008 = \in185  & n1787;
  assign n2009 = \in085  & ~n1787;
  assign n2010 = ~n2008 & ~n2009;
  assign n2011 = \in385  & n1792;
  assign n2012 = \in285  & ~n1792;
  assign n2013 = ~n2011 & ~n2012;
  assign n2014 = n2010 & ~n2013;
  assign n2015 = \in184  & n1787;
  assign n2016 = \in084  & ~n1787;
  assign n2017 = ~n2015 & ~n2016;
  assign n2018 = \in384  & n1792;
  assign n2019 = \in284  & ~n1792;
  assign n2020 = ~n2018 & ~n2019;
  assign n2021 = ~n2017 & n2020;
  assign n2022 = ~n2014 & n2021;
  assign n2023 = ~n2010 & n2013;
  assign n2024 = ~n2022 & ~n2023;
  assign n2025 = n2007 & ~n2024;
  assign n2026 = n2002 & ~n2005;
  assign n2027 = ~n1999 & n2026;
  assign n2028 = \in380  & n1792;
  assign n2029 = \in280  & ~n1792;
  assign n2030 = ~n2028 & ~n2029;
  assign n2031 = \in180  & n1787;
  assign n2032 = \in080  & ~n1787;
  assign n2033 = ~n2031 & ~n2032;
  assign n2034 = ~n2030 & n2033;
  assign n2035 = \in183  & n1787;
  assign n2036 = \in083  & ~n1787;
  assign n2037 = ~n2035 & ~n2036;
  assign n2038 = \in383  & n1792;
  assign n2039 = \in283  & ~n1792;
  assign n2040 = ~n2038 & ~n2039;
  assign n2041 = n2037 & ~n2040;
  assign n2042 = \in382  & n1792;
  assign n2043 = \in282  & ~n1792;
  assign n2044 = ~n2042 & ~n2043;
  assign n2045 = \in182  & n1787;
  assign n2046 = \in082  & ~n1787;
  assign n2047 = ~n2045 & ~n2046;
  assign n2048 = ~n2044 & n2047;
  assign n2049 = ~n2041 & ~n2048;
  assign n2050 = \in181  & n1787;
  assign n2051 = \in081  & ~n1787;
  assign n2052 = ~n2050 & ~n2051;
  assign n2053 = \in381  & n1792;
  assign n2054 = \in281  & ~n1792;
  assign n2055 = ~n2053 & ~n2054;
  assign n2056 = n2052 & ~n2055;
  assign n2057 = \in179  & n1787;
  assign n2058 = \in079  & ~n1787;
  assign n2059 = ~n2057 & ~n2058;
  assign n2060 = \in379  & n1792;
  assign n2061 = \in279  & ~n1792;
  assign n2062 = ~n2060 & ~n2061;
  assign n2063 = ~n2059 & n2062;
  assign n2064 = n2059 & ~n2062;
  assign n2065 = \in378  & n1792;
  assign n2066 = \in278  & ~n1792;
  assign n2067 = ~n2065 & ~n2066;
  assign n2068 = \in178  & n1787;
  assign n2069 = \in078  & ~n1787;
  assign n2070 = ~n2068 & ~n2069;
  assign n2071 = ~n2067 & n2070;
  assign n2072 = ~n2064 & ~n2071;
  assign n2073 = \in177  & n1787;
  assign n2074 = \in077  & ~n1787;
  assign n2075 = ~n2073 & ~n2074;
  assign n2076 = \in377  & n1792;
  assign n2077 = \in277  & ~n1792;
  assign n2078 = ~n2076 & ~n2077;
  assign n2079 = n2075 & ~n2078;
  assign n2080 = \in176  & n1787;
  assign n2081 = \in076  & ~n1787;
  assign n2082 = ~n2080 & ~n2081;
  assign n2083 = \in376  & n1792;
  assign n2084 = \in276  & ~n1792;
  assign n2085 = ~n2083 & ~n2084;
  assign n2086 = ~n2082 & n2085;
  assign n2087 = ~n2079 & n2086;
  assign n2088 = ~n2075 & n2078;
  assign n2089 = ~n2087 & ~n2088;
  assign n2090 = n2072 & ~n2089;
  assign n2091 = n2067 & ~n2070;
  assign n2092 = ~n2064 & n2091;
  assign n2093 = \in171  & n1787;
  assign n2094 = \in071  & ~n1787;
  assign n2095 = ~n2093 & ~n2094;
  assign n2096 = \in371  & n1792;
  assign n2097 = \in271  & ~n1792;
  assign n2098 = ~n2096 & ~n2097;
  assign n2099 = ~n2095 & n2098;
  assign n2100 = n2095 & ~n2098;
  assign n2101 = \in370  & n1792;
  assign n2102 = \in270  & ~n1792;
  assign n2103 = ~n2101 & ~n2102;
  assign n2104 = \in170  & n1787;
  assign n2105 = \in070  & ~n1787;
  assign n2106 = ~n2104 & ~n2105;
  assign n2107 = ~n2103 & n2106;
  assign n2108 = ~n2100 & ~n2107;
  assign n2109 = \in169  & n1787;
  assign n2110 = \in069  & ~n1787;
  assign n2111 = ~n2109 & ~n2110;
  assign n2112 = \in369  & n1792;
  assign n2113 = \in269  & ~n1792;
  assign n2114 = ~n2112 & ~n2113;
  assign n2115 = n2111 & ~n2114;
  assign n2116 = \in168  & n1787;
  assign n2117 = \in068  & ~n1787;
  assign n2118 = ~n2116 & ~n2117;
  assign n2119 = \in368  & n1792;
  assign n2120 = \in268  & ~n1792;
  assign n2121 = ~n2119 & ~n2120;
  assign n2122 = ~n2118 & n2121;
  assign n2123 = ~n2115 & n2122;
  assign n2124 = ~n2111 & n2114;
  assign n2125 = ~n2123 & ~n2124;
  assign n2126 = n2108 & ~n2125;
  assign n2127 = n2103 & ~n2106;
  assign n2128 = ~n2100 & n2127;
  assign n2129 = \in167  & n1787;
  assign n2130 = \in067  & ~n1787;
  assign n2131 = ~n2129 & ~n2130;
  assign n2132 = \in367  & n1792;
  assign n2133 = \in267  & ~n1792;
  assign n2134 = ~n2132 & ~n2133;
  assign n2135 = n2131 & ~n2134;
  assign n2136 = \in366  & n1792;
  assign n2137 = \in266  & ~n1792;
  assign n2138 = ~n2136 & ~n2137;
  assign n2139 = \in166  & n1787;
  assign n2140 = \in066  & ~n1787;
  assign n2141 = ~n2139 & ~n2140;
  assign n2142 = ~n2138 & n2141;
  assign n2143 = ~n2135 & ~n2142;
  assign n2144 = \in364  & n1792;
  assign n2145 = \in264  & ~n1792;
  assign n2146 = ~n2144 & ~n2145;
  assign n2147 = \in164  & n1787;
  assign n2148 = \in064  & ~n1787;
  assign n2149 = ~n2147 & ~n2148;
  assign n2150 = ~n2146 & n2149;
  assign n2151 = \in165  & n1787;
  assign n2152 = \in065  & ~n1787;
  assign n2153 = ~n2151 & ~n2152;
  assign n2154 = \in365  & n1792;
  assign n2155 = \in265  & ~n1792;
  assign n2156 = ~n2154 & ~n2155;
  assign n2157 = n2153 & ~n2156;
  assign n2158 = \in163  & n1787;
  assign n2159 = \in063  & ~n1787;
  assign n2160 = ~n2158 & ~n2159;
  assign n2161 = \in363  & n1792;
  assign n2162 = \in263  & ~n1792;
  assign n2163 = ~n2161 & ~n2162;
  assign n2164 = ~n2160 & n2163;
  assign n2165 = n2160 & ~n2163;
  assign n2166 = \in362  & n1792;
  assign n2167 = \in262  & ~n1792;
  assign n2168 = ~n2166 & ~n2167;
  assign n2169 = \in162  & n1787;
  assign n2170 = \in062  & ~n1787;
  assign n2171 = ~n2169 & ~n2170;
  assign n2172 = ~n2168 & n2171;
  assign n2173 = ~n2165 & ~n2172;
  assign n2174 = \in160  & n1787;
  assign n2175 = \in060  & ~n1787;
  assign n2176 = ~n2174 & ~n2175;
  assign n2177 = \in360  & n1792;
  assign n2178 = \in260  & ~n1792;
  assign n2179 = ~n2177 & ~n2178;
  assign n2180 = n2176 & ~n2179;
  assign n2181 = \in161  & n1787;
  assign n2182 = \in061  & ~n1787;
  assign n2183 = ~n2181 & ~n2182;
  assign n2184 = \in361  & n1792;
  assign n2185 = \in261  & ~n1792;
  assign n2186 = ~n2184 & ~n2185;
  assign n2187 = n2183 & ~n2186;
  assign n2188 = ~n2180 & ~n2187;
  assign n2189 = n2173 & n2188;
  assign n2190 = \in159  & n1787;
  assign n2191 = \in059  & ~n1787;
  assign n2192 = ~n2190 & ~n2191;
  assign n2193 = \in359  & n1792;
  assign n2194 = \in259  & ~n1792;
  assign n2195 = ~n2193 & ~n2194;
  assign n2196 = ~n2192 & n2195;
  assign n2197 = n2192 & ~n2195;
  assign n2198 = \in158  & n1787;
  assign n2199 = \in058  & ~n1787;
  assign n2200 = ~n2198 & ~n2199;
  assign n2201 = \in358  & n1792;
  assign n2202 = \in258  & ~n1792;
  assign n2203 = ~n2201 & ~n2202;
  assign n2204 = n2200 & ~n2203;
  assign n2205 = ~n2197 & ~n2204;
  assign n2206 = \in157  & n1787;
  assign n2207 = \in057  & ~n1787;
  assign n2208 = ~n2206 & ~n2207;
  assign n2209 = \in357  & n1792;
  assign n2210 = \in257  & ~n1792;
  assign n2211 = ~n2209 & ~n2210;
  assign n2212 = n2208 & ~n2211;
  assign n2213 = \in156  & n1787;
  assign n2214 = \in056  & ~n1787;
  assign n2215 = ~n2213 & ~n2214;
  assign n2216 = \in356  & n1792;
  assign n2217 = \in256  & ~n1792;
  assign n2218 = ~n2216 & ~n2217;
  assign n2219 = ~n2215 & n2218;
  assign n2220 = ~n2212 & n2219;
  assign n2221 = ~n2208 & n2211;
  assign n2222 = ~n2220 & ~n2221;
  assign n2223 = ~n2200 & n2203;
  assign n2224 = n2222 & ~n2223;
  assign n2225 = n2205 & ~n2224;
  assign n2226 = ~n2196 & ~n2225;
  assign n2227 = n2189 & ~n2226;
  assign n2228 = ~n2176 & n2179;
  assign n2229 = ~n2187 & n2228;
  assign n2230 = ~n2183 & n2186;
  assign n2231 = ~n2229 & ~n2230;
  assign n2232 = n2173 & ~n2231;
  assign n2233 = n2168 & ~n2171;
  assign n2234 = ~n2165 & n2233;
  assign n2235 = \in147  & n1787;
  assign n2236 = \in047  & ~n1787;
  assign n2237 = ~n2235 & ~n2236;
  assign n2238 = \in347  & n1792;
  assign n2239 = \in247  & ~n1792;
  assign n2240 = ~n2238 & ~n2239;
  assign n2241 = ~n2237 & n2240;
  assign n2242 = n2237 & ~n2240;
  assign n2243 = \in346  & n1792;
  assign n2244 = \in246  & ~n1792;
  assign n2245 = ~n2243 & ~n2244;
  assign n2246 = \in146  & n1787;
  assign n2247 = \in046  & ~n1787;
  assign n2248 = ~n2246 & ~n2247;
  assign n2249 = ~n2245 & n2248;
  assign n2250 = ~n2242 & ~n2249;
  assign n2251 = \in144  & n1787;
  assign n2252 = \in044  & ~n1787;
  assign n2253 = ~n2251 & ~n2252;
  assign n2254 = \in344  & n1792;
  assign n2255 = \in244  & ~n1792;
  assign n2256 = ~n2254 & ~n2255;
  assign n2257 = n2253 & ~n2256;
  assign n2258 = \in145  & n1787;
  assign n2259 = \in045  & ~n1787;
  assign n2260 = ~n2258 & ~n2259;
  assign n2261 = \in345  & n1792;
  assign n2262 = \in245  & ~n1792;
  assign n2263 = ~n2261 & ~n2262;
  assign n2264 = n2260 & ~n2263;
  assign n2265 = ~n2257 & ~n2264;
  assign n2266 = n2250 & n2265;
  assign n2267 = \in143  & n1787;
  assign n2268 = \in043  & ~n1787;
  assign n2269 = ~n2267 & ~n2268;
  assign n2270 = \in343  & n1792;
  assign n2271 = \in243  & ~n1792;
  assign n2272 = ~n2270 & ~n2271;
  assign n2273 = ~n2269 & n2272;
  assign n2274 = n2269 & ~n2272;
  assign n2275 = \in142  & n1787;
  assign n2276 = \in042  & ~n1787;
  assign n2277 = ~n2275 & ~n2276;
  assign n2278 = \in342  & n1792;
  assign n2279 = \in242  & ~n1792;
  assign n2280 = ~n2278 & ~n2279;
  assign n2281 = n2277 & ~n2280;
  assign n2282 = ~n2274 & ~n2281;
  assign n2283 = \in141  & n1787;
  assign n2284 = \in041  & ~n1787;
  assign n2285 = ~n2283 & ~n2284;
  assign n2286 = \in341  & n1792;
  assign n2287 = \in241  & ~n1792;
  assign n2288 = ~n2286 & ~n2287;
  assign n2289 = n2285 & ~n2288;
  assign n2290 = \in140  & n1787;
  assign n2291 = \in040  & ~n1787;
  assign n2292 = ~n2290 & ~n2291;
  assign n2293 = \in340  & n1792;
  assign n2294 = \in240  & ~n1792;
  assign n2295 = ~n2293 & ~n2294;
  assign n2296 = ~n2292 & n2295;
  assign n2297 = ~n2289 & n2296;
  assign n2298 = ~n2285 & n2288;
  assign n2299 = ~n2297 & ~n2298;
  assign n2300 = ~n2277 & n2280;
  assign n2301 = n2299 & ~n2300;
  assign n2302 = n2282 & ~n2301;
  assign n2303 = ~n2273 & ~n2302;
  assign n2304 = n2266 & ~n2303;
  assign n2305 = ~n2253 & n2256;
  assign n2306 = ~n2264 & n2305;
  assign n2307 = ~n2260 & n2263;
  assign n2308 = ~n2306 & ~n2307;
  assign n2309 = n2250 & ~n2308;
  assign n2310 = n2245 & ~n2248;
  assign n2311 = ~n2242 & n2310;
  assign n2312 = \in332  & n1792;
  assign n2313 = \in232  & ~n1792;
  assign n2314 = ~n2312 & ~n2313;
  assign n2315 = \in132  & n1787;
  assign n2316 = \in032  & ~n1787;
  assign n2317 = ~n2315 & ~n2316;
  assign n2318 = ~n2314 & n2317;
  assign n2319 = \in131  & n1787;
  assign n2320 = \in031  & ~n1787;
  assign n2321 = ~n2319 & ~n2320;
  assign n2322 = \in331  & n1792;
  assign n2323 = \in231  & ~n1792;
  assign n2324 = ~n2322 & ~n2323;
  assign n2325 = n2321 & ~n2324;
  assign n2326 = \in130  & n1787;
  assign n2327 = \in030  & ~n1787;
  assign n2328 = ~n2326 & ~n2327;
  assign n2329 = \in330  & n1792;
  assign n2330 = \in230  & ~n1792;
  assign n2331 = ~n2329 & ~n2330;
  assign n2332 = n2328 & ~n2331;
  assign n2333 = \in129  & n1787;
  assign n2334 = \in029  & ~n1787;
  assign n2335 = ~n2333 & ~n2334;
  assign n2336 = \in329  & n1792;
  assign n2337 = \in229  & ~n1792;
  assign n2338 = ~n2336 & ~n2337;
  assign n2339 = n2335 & ~n2338;
  assign n2340 = \in128  & n1787;
  assign n2341 = \in028  & ~n1787;
  assign n2342 = ~n2340 & ~n2341;
  assign n2343 = \in328  & n1792;
  assign n2344 = \in228  & ~n1792;
  assign n2345 = ~n2343 & ~n2344;
  assign n2346 = n2342 & ~n2345;
  assign n2347 = \in127  & n1787;
  assign n2348 = \in027  & ~n1787;
  assign n2349 = ~n2347 & ~n2348;
  assign n2350 = \in327  & n1792;
  assign n2351 = \in227  & ~n1792;
  assign n2352 = ~n2350 & ~n2351;
  assign n2353 = n2349 & ~n2352;
  assign n2354 = \in126  & n1787;
  assign n2355 = \in026  & ~n1787;
  assign n2356 = ~n2354 & ~n2355;
  assign n2357 = \in326  & n1792;
  assign n2358 = \in226  & ~n1792;
  assign n2359 = ~n2357 & ~n2358;
  assign n2360 = n2356 & ~n2359;
  assign n2361 = \in325  & n1792;
  assign n2362 = \in225  & ~n1792;
  assign n2363 = ~n2361 & ~n2362;
  assign n2364 = \in324  & n1792;
  assign n2365 = \in224  & ~n1792;
  assign n2366 = ~n2364 & ~n2365;
  assign n2367 = \in123  & n1787;
  assign n2368 = \in023  & ~n1787;
  assign n2369 = ~n2367 & ~n2368;
  assign n2370 = \in323  & n1792;
  assign n2371 = \in223  & ~n1792;
  assign n2372 = ~n2370 & ~n2371;
  assign n2373 = n2369 & ~n2372;
  assign n2374 = \in122  & n1787;
  assign n2375 = \in022  & ~n1787;
  assign n2376 = ~n2374 & ~n2375;
  assign n2377 = \in322  & n1792;
  assign n2378 = \in222  & ~n1792;
  assign n2379 = ~n2377 & ~n2378;
  assign n2380 = n2376 & ~n2379;
  assign n2381 = \in121  & n1787;
  assign n2382 = \in021  & ~n1787;
  assign n2383 = ~n2381 & ~n2382;
  assign n2384 = \in321  & n1792;
  assign n2385 = \in221  & ~n1792;
  assign n2386 = ~n2384 & ~n2385;
  assign n2387 = n2383 & ~n2386;
  assign n2388 = \in120  & n1787;
  assign n2389 = \in020  & ~n1787;
  assign n2390 = ~n2388 & ~n2389;
  assign n2391 = \in320  & n1792;
  assign n2392 = \in220  & ~n1792;
  assign n2393 = ~n2391 & ~n2392;
  assign n2394 = n2390 & ~n2393;
  assign n2395 = \in119  & n1787;
  assign n2396 = \in019  & ~n1787;
  assign n2397 = ~n2395 & ~n2396;
  assign n2398 = \in319  & n1792;
  assign n2399 = \in219  & ~n1792;
  assign n2400 = ~n2398 & ~n2399;
  assign n2401 = n2397 & ~n2400;
  assign n2402 = \in118  & n1787;
  assign n2403 = \in018  & ~n1787;
  assign n2404 = ~n2402 & ~n2403;
  assign n2405 = \in318  & n1792;
  assign n2406 = \in218  & ~n1792;
  assign n2407 = ~n2405 & ~n2406;
  assign n2408 = n2404 & ~n2407;
  assign n2409 = \in317  & n1792;
  assign n2410 = \in217  & ~n1792;
  assign n2411 = ~n2409 & ~n2410;
  assign n2412 = \in316  & n1792;
  assign n2413 = \in216  & ~n1792;
  assign n2414 = ~n2412 & ~n2413;
  assign n2415 = \in115  & n1787;
  assign n2416 = \in015  & ~n1787;
  assign n2417 = ~n2415 & ~n2416;
  assign n2418 = \in315  & n1792;
  assign n2419 = \in215  & ~n1792;
  assign n2420 = ~n2418 & ~n2419;
  assign n2421 = n2417 & ~n2420;
  assign n2422 = \in114  & n1787;
  assign n2423 = \in014  & ~n1787;
  assign n2424 = ~n2422 & ~n2423;
  assign n2425 = \in314  & n1792;
  assign n2426 = \in214  & ~n1792;
  assign n2427 = ~n2425 & ~n2426;
  assign n2428 = n2424 & ~n2427;
  assign n2429 = \in113  & n1787;
  assign n2430 = \in013  & ~n1787;
  assign n2431 = ~n2429 & ~n2430;
  assign n2432 = \in313  & n1792;
  assign n2433 = \in213  & ~n1792;
  assign n2434 = ~n2432 & ~n2433;
  assign n2435 = n2431 & ~n2434;
  assign n2436 = \in112  & n1787;
  assign n2437 = \in012  & ~n1787;
  assign n2438 = ~n2436 & ~n2437;
  assign n2439 = \in312  & n1792;
  assign n2440 = \in212  & ~n1792;
  assign n2441 = ~n2439 & ~n2440;
  assign n2442 = n2438 & ~n2441;
  assign n2443 = \in111  & n1787;
  assign n2444 = \in011  & ~n1787;
  assign n2445 = ~n2443 & ~n2444;
  assign n2446 = \in311  & n1792;
  assign n2447 = \in211  & ~n1792;
  assign n2448 = ~n2446 & ~n2447;
  assign n2449 = n2445 & ~n2448;
  assign n2450 = \in110  & n1787;
  assign n2451 = \in010  & ~n1787;
  assign n2452 = ~n2450 & ~n2451;
  assign n2453 = \in310  & n1792;
  assign n2454 = \in210  & ~n1792;
  assign n2455 = ~n2453 & ~n2454;
  assign n2456 = n2452 & ~n2455;
  assign n2457 = \in39  & n1792;
  assign n2458 = \in29  & ~n1792;
  assign n2459 = ~n2457 & ~n2458;
  assign n2460 = \in38  & n1792;
  assign n2461 = \in28  & ~n1792;
  assign n2462 = ~n2460 & ~n2461;
  assign n2463 = \in17  & n1787;
  assign n2464 = \in07  & ~n1787;
  assign n2465 = ~n2463 & ~n2464;
  assign n2466 = \in37  & n1792;
  assign n2467 = \in27  & ~n1792;
  assign n2468 = ~n2466 & ~n2467;
  assign n2469 = n2465 & ~n2468;
  assign n2470 = \in36  & n1792;
  assign n2471 = \in26  & ~n1792;
  assign n2472 = ~n2470 & ~n2471;
  assign n2473 = \in16  & n1787;
  assign n2474 = \in06  & ~n1787;
  assign n2475 = ~n2473 & ~n2474;
  assign n2476 = \in35  & n1792;
  assign n2477 = \in25  & ~n1792;
  assign n2478 = ~n2476 & ~n2477;
  assign n2479 = \in15  & n1787;
  assign n2480 = \in05  & ~n1787;
  assign n2481 = ~n2479 & ~n2480;
  assign n2482 = \in34  & n1792;
  assign n2483 = \in24  & ~n1792;
  assign n2484 = ~n2482 & ~n2483;
  assign n2485 = \in14  & n1787;
  assign n2486 = \in04  & ~n1787;
  assign n2487 = ~n2485 & ~n2486;
  assign n2488 = \in13  & n1787;
  assign n2489 = \in03  & ~n1787;
  assign n2490 = ~n2488 & ~n2489;
  assign n2491 = \in33  & n1792;
  assign n2492 = \in23  & ~n1792;
  assign n2493 = ~n2491 & ~n2492;
  assign n2494 = n2490 & ~n2493;
  assign n2495 = \in31  & n1792;
  assign n2496 = \in21  & ~n1792;
  assign n2497 = ~n2495 & ~n2496;
  assign n2498 = \in10  & n1787;
  assign n2499 = \in00  & ~n1787;
  assign n2500 = ~n2498 & ~n2499;
  assign n2501 = \in30  & n1792;
  assign n2502 = \in20  & ~n1792;
  assign n2503 = ~n2501 & ~n2502;
  assign n2504 = ~n2500 & n2503;
  assign n2505 = n2497 & n2504;
  assign n2506 = \in11  & n1787;
  assign n2507 = \in01  & ~n1787;
  assign n2508 = ~n2506 & ~n2507;
  assign n2509 = ~n2505 & n2508;
  assign n2510 = \in12  & n1787;
  assign n2511 = \in02  & ~n1787;
  assign n2512 = ~n2510 & ~n2511;
  assign n2513 = \in32  & n1792;
  assign n2514 = \in22  & ~n1792;
  assign n2515 = ~n2513 & ~n2514;
  assign n2516 = n2512 & ~n2515;
  assign n2517 = ~n2497 & ~n2504;
  assign n2518 = ~n2516 & ~n2517;
  assign n2519 = ~n2509 & n2518;
  assign n2520 = ~n2512 & n2515;
  assign n2521 = ~n2519 & ~n2520;
  assign n2522 = ~n2494 & ~n2521;
  assign n2523 = ~n2490 & n2493;
  assign n2524 = ~n2522 & ~n2523;
  assign n2525 = n2487 & n2524;
  assign n2526 = n2484 & ~n2525;
  assign n2527 = ~n2487 & ~n2524;
  assign n2528 = ~n2526 & ~n2527;
  assign n2529 = n2481 & n2528;
  assign n2530 = n2478 & ~n2529;
  assign n2531 = ~n2481 & ~n2528;
  assign n2532 = ~n2530 & ~n2531;
  assign n2533 = n2475 & n2532;
  assign n2534 = n2472 & ~n2533;
  assign n2535 = ~n2475 & ~n2532;
  assign n2536 = ~n2534 & ~n2535;
  assign n2537 = ~n2469 & ~n2536;
  assign n2538 = ~n2465 & n2468;
  assign n2539 = ~n2537 & ~n2538;
  assign n2540 = \in18  & n1787;
  assign n2541 = \in08  & ~n1787;
  assign n2542 = ~n2540 & ~n2541;
  assign n2543 = n2539 & n2542;
  assign n2544 = n2462 & ~n2543;
  assign n2545 = ~n2539 & ~n2542;
  assign n2546 = ~n2544 & ~n2545;
  assign n2547 = \in19  & n1787;
  assign n2548 = \in09  & ~n1787;
  assign n2549 = ~n2547 & ~n2548;
  assign n2550 = n2546 & n2549;
  assign n2551 = n2459 & ~n2550;
  assign n2552 = ~n2546 & ~n2549;
  assign n2553 = ~n2551 & ~n2552;
  assign n2554 = ~n2456 & ~n2553;
  assign n2555 = ~n2452 & n2455;
  assign n2556 = ~n2554 & ~n2555;
  assign n2557 = ~n2449 & ~n2556;
  assign n2558 = ~n2445 & n2448;
  assign n2559 = ~n2557 & ~n2558;
  assign n2560 = ~n2442 & ~n2559;
  assign n2561 = ~n2438 & n2441;
  assign n2562 = ~n2560 & ~n2561;
  assign n2563 = ~n2435 & ~n2562;
  assign n2564 = ~n2431 & n2434;
  assign n2565 = ~n2563 & ~n2564;
  assign n2566 = ~n2428 & ~n2565;
  assign n2567 = ~n2424 & n2427;
  assign n2568 = ~n2566 & ~n2567;
  assign n2569 = ~n2421 & ~n2568;
  assign n2570 = ~n2417 & n2420;
  assign n2571 = ~n2569 & ~n2570;
  assign n2572 = \in116  & n1787;
  assign n2573 = \in016  & ~n1787;
  assign n2574 = ~n2572 & ~n2573;
  assign n2575 = n2571 & n2574;
  assign n2576 = n2414 & ~n2575;
  assign n2577 = ~n2571 & ~n2574;
  assign n2578 = ~n2576 & ~n2577;
  assign n2579 = \in117  & n1787;
  assign n2580 = \in017  & ~n1787;
  assign n2581 = ~n2579 & ~n2580;
  assign n2582 = n2578 & n2581;
  assign n2583 = n2411 & ~n2582;
  assign n2584 = ~n2578 & ~n2581;
  assign n2585 = ~n2583 & ~n2584;
  assign n2586 = ~n2408 & ~n2585;
  assign n2587 = ~n2404 & n2407;
  assign n2588 = ~n2586 & ~n2587;
  assign n2589 = ~n2401 & ~n2588;
  assign n2590 = ~n2397 & n2400;
  assign n2591 = ~n2589 & ~n2590;
  assign n2592 = ~n2394 & ~n2591;
  assign n2593 = ~n2390 & n2393;
  assign n2594 = ~n2592 & ~n2593;
  assign n2595 = ~n2387 & ~n2594;
  assign n2596 = ~n2383 & n2386;
  assign n2597 = ~n2595 & ~n2596;
  assign n2598 = ~n2380 & ~n2597;
  assign n2599 = ~n2376 & n2379;
  assign n2600 = ~n2598 & ~n2599;
  assign n2601 = ~n2373 & ~n2600;
  assign n2602 = ~n2369 & n2372;
  assign n2603 = ~n2601 & ~n2602;
  assign n2604 = \in124  & n1787;
  assign n2605 = \in024  & ~n1787;
  assign n2606 = ~n2604 & ~n2605;
  assign n2607 = n2603 & n2606;
  assign n2608 = n2366 & ~n2607;
  assign n2609 = ~n2603 & ~n2606;
  assign n2610 = ~n2608 & ~n2609;
  assign n2611 = \in125  & n1787;
  assign n2612 = \in025  & ~n1787;
  assign n2613 = ~n2611 & ~n2612;
  assign n2614 = n2610 & n2613;
  assign n2615 = n2363 & ~n2614;
  assign n2616 = ~n2610 & ~n2613;
  assign n2617 = ~n2615 & ~n2616;
  assign n2618 = ~n2360 & ~n2617;
  assign n2619 = ~n2356 & n2359;
  assign n2620 = ~n2618 & ~n2619;
  assign n2621 = ~n2353 & ~n2620;
  assign n2622 = ~n2349 & n2352;
  assign n2623 = ~n2621 & ~n2622;
  assign n2624 = ~n2346 & ~n2623;
  assign n2625 = ~n2342 & n2345;
  assign n2626 = ~n2624 & ~n2625;
  assign n2627 = ~n2339 & ~n2626;
  assign n2628 = ~n2335 & n2338;
  assign n2629 = ~n2627 & ~n2628;
  assign n2630 = ~n2332 & ~n2629;
  assign n2631 = ~n2328 & n2331;
  assign n2632 = ~n2630 & ~n2631;
  assign n2633 = ~n2325 & ~n2632;
  assign n2634 = ~n2321 & n2324;
  assign n2635 = ~n2633 & ~n2634;
  assign n2636 = \in139  & n1787;
  assign n2637 = \in039  & ~n1787;
  assign n2638 = ~n2636 & ~n2637;
  assign n2639 = \in339  & n1792;
  assign n2640 = \in239  & ~n1792;
  assign n2641 = ~n2639 & ~n2640;
  assign n2642 = n2638 & ~n2641;
  assign n2643 = \in338  & n1792;
  assign n2644 = \in238  & ~n1792;
  assign n2645 = ~n2643 & ~n2644;
  assign n2646 = \in138  & n1787;
  assign n2647 = \in038  & ~n1787;
  assign n2648 = ~n2646 & ~n2647;
  assign n2649 = ~n2645 & n2648;
  assign n2650 = ~n2642 & ~n2649;
  assign n2651 = \in136  & n1787;
  assign n2652 = \in036  & ~n1787;
  assign n2653 = ~n2651 & ~n2652;
  assign n2654 = \in336  & n1792;
  assign n2655 = \in236  & ~n1792;
  assign n2656 = ~n2654 & ~n2655;
  assign n2657 = n2653 & ~n2656;
  assign n2658 = \in137  & n1787;
  assign n2659 = \in037  & ~n1787;
  assign n2660 = ~n2658 & ~n2659;
  assign n2661 = \in337  & n1792;
  assign n2662 = \in237  & ~n1792;
  assign n2663 = ~n2661 & ~n2662;
  assign n2664 = n2660 & ~n2663;
  assign n2665 = ~n2657 & ~n2664;
  assign n2666 = n2650 & n2665;
  assign n2667 = \in133  & n1787;
  assign n2668 = \in033  & ~n1787;
  assign n2669 = ~n2667 & ~n2668;
  assign n2670 = \in333  & n1792;
  assign n2671 = \in233  & ~n1792;
  assign n2672 = ~n2670 & ~n2671;
  assign n2673 = n2669 & ~n2672;
  assign n2674 = \in135  & n1787;
  assign n2675 = \in035  & ~n1787;
  assign n2676 = ~n2674 & ~n2675;
  assign n2677 = \in335  & n1792;
  assign n2678 = \in235  & ~n1792;
  assign n2679 = ~n2677 & ~n2678;
  assign n2680 = n2676 & ~n2679;
  assign n2681 = \in334  & n1792;
  assign n2682 = \in234  & ~n1792;
  assign n2683 = ~n2681 & ~n2682;
  assign n2684 = \in134  & n1787;
  assign n2685 = \in034  & ~n1787;
  assign n2686 = ~n2684 & ~n2685;
  assign n2687 = ~n2683 & n2686;
  assign n2688 = ~n2680 & ~n2687;
  assign n2689 = ~n2673 & n2688;
  assign n2690 = n2666 & n2689;
  assign n2691 = ~n2635 & n2690;
  assign n2692 = ~n2318 & n2691;
  assign n2693 = ~n2638 & n2641;
  assign n2694 = ~n2653 & n2656;
  assign n2695 = ~n2664 & n2694;
  assign n2696 = ~n2660 & n2663;
  assign n2697 = ~n2695 & ~n2696;
  assign n2698 = n2650 & ~n2697;
  assign n2699 = ~n2642 & n2645;
  assign n2700 = ~n2648 & n2699;
  assign n2701 = ~n2676 & n2679;
  assign n2702 = ~n2680 & n2683;
  assign n2703 = ~n2686 & n2702;
  assign n2704 = n2314 & ~n2317;
  assign n2705 = ~n2669 & n2672;
  assign n2706 = ~n2704 & ~n2705;
  assign n2707 = n2689 & ~n2706;
  assign n2708 = ~n2703 & ~n2707;
  assign n2709 = ~n2701 & n2708;
  assign n2710 = n2666 & ~n2709;
  assign n2711 = ~n2700 & ~n2710;
  assign n2712 = ~n2698 & n2711;
  assign n2713 = ~n2693 & n2712;
  assign n2714 = ~n2692 & n2713;
  assign n2715 = n2292 & ~n2295;
  assign n2716 = ~n2289 & ~n2715;
  assign n2717 = n2282 & n2716;
  assign n2718 = n2266 & n2717;
  assign n2719 = ~n2714 & n2718;
  assign n2720 = ~n2311 & ~n2719;
  assign n2721 = ~n2309 & n2720;
  assign n2722 = ~n2304 & n2721;
  assign n2723 = ~n2241 & n2722;
  assign n2724 = \in348  & n1792;
  assign n2725 = \in248  & ~n1792;
  assign n2726 = ~n2724 & ~n2725;
  assign n2727 = \in148  & n1787;
  assign n2728 = \in048  & ~n1787;
  assign n2729 = ~n2727 & ~n2728;
  assign n2730 = ~n2726 & n2729;
  assign n2731 = \in155  & n1787;
  assign n2732 = \in055  & ~n1787;
  assign n2733 = ~n2731 & ~n2732;
  assign n2734 = \in355  & n1792;
  assign n2735 = \in255  & ~n1792;
  assign n2736 = ~n2734 & ~n2735;
  assign n2737 = n2733 & ~n2736;
  assign n2738 = \in354  & n1792;
  assign n2739 = \in254  & ~n1792;
  assign n2740 = ~n2738 & ~n2739;
  assign n2741 = \in154  & n1787;
  assign n2742 = \in054  & ~n1787;
  assign n2743 = ~n2741 & ~n2742;
  assign n2744 = ~n2740 & n2743;
  assign n2745 = ~n2737 & ~n2744;
  assign n2746 = \in153  & n1787;
  assign n2747 = \in053  & ~n1787;
  assign n2748 = ~n2746 & ~n2747;
  assign n2749 = \in353  & n1792;
  assign n2750 = \in253  & ~n1792;
  assign n2751 = ~n2749 & ~n2750;
  assign n2752 = n2748 & ~n2751;
  assign n2753 = \in352  & n1792;
  assign n2754 = \in252  & ~n1792;
  assign n2755 = ~n2753 & ~n2754;
  assign n2756 = \in152  & n1787;
  assign n2757 = \in052  & ~n1787;
  assign n2758 = ~n2756 & ~n2757;
  assign n2759 = ~n2755 & n2758;
  assign n2760 = ~n2752 & ~n2759;
  assign n2761 = n2745 & n2760;
  assign n2762 = \in149  & n1787;
  assign n2763 = \in049  & ~n1787;
  assign n2764 = ~n2762 & ~n2763;
  assign n2765 = \in349  & n1792;
  assign n2766 = \in249  & ~n1792;
  assign n2767 = ~n2765 & ~n2766;
  assign n2768 = n2764 & ~n2767;
  assign n2769 = \in151  & n1787;
  assign n2770 = \in051  & ~n1787;
  assign n2771 = ~n2769 & ~n2770;
  assign n2772 = \in351  & n1792;
  assign n2773 = \in251  & ~n1792;
  assign n2774 = ~n2772 & ~n2773;
  assign n2775 = n2771 & ~n2774;
  assign n2776 = \in350  & n1792;
  assign n2777 = \in250  & ~n1792;
  assign n2778 = ~n2776 & ~n2777;
  assign n2779 = \in150  & n1787;
  assign n2780 = \in050  & ~n1787;
  assign n2781 = ~n2779 & ~n2780;
  assign n2782 = ~n2778 & n2781;
  assign n2783 = ~n2775 & ~n2782;
  assign n2784 = ~n2768 & n2783;
  assign n2785 = n2761 & n2784;
  assign n2786 = ~n2730 & n2785;
  assign n2787 = ~n2723 & n2786;
  assign n2788 = ~n2733 & n2736;
  assign n2789 = ~n2771 & n2774;
  assign n2790 = ~n2775 & n2778;
  assign n2791 = ~n2781 & n2790;
  assign n2792 = n2726 & ~n2729;
  assign n2793 = ~n2764 & n2767;
  assign n2794 = ~n2792 & ~n2793;
  assign n2795 = n2784 & ~n2794;
  assign n2796 = ~n2791 & ~n2795;
  assign n2797 = ~n2789 & n2796;
  assign n2798 = n2761 & ~n2797;
  assign n2799 = n2755 & ~n2758;
  assign n2800 = ~n2752 & n2799;
  assign n2801 = ~n2748 & n2751;
  assign n2802 = ~n2800 & ~n2801;
  assign n2803 = n2740 & ~n2743;
  assign n2804 = n2802 & ~n2803;
  assign n2805 = n2745 & ~n2804;
  assign n2806 = ~n2798 & ~n2805;
  assign n2807 = ~n2788 & n2806;
  assign n2808 = ~n2787 & n2807;
  assign n2809 = n2215 & ~n2218;
  assign n2810 = ~n2212 & ~n2809;
  assign n2811 = n2189 & n2810;
  assign n2812 = n2205 & n2811;
  assign n2813 = ~n2808 & n2812;
  assign n2814 = ~n2234 & ~n2813;
  assign n2815 = ~n2232 & n2814;
  assign n2816 = ~n2227 & n2815;
  assign n2817 = ~n2164 & n2816;
  assign n2818 = ~n2157 & ~n2817;
  assign n2819 = ~n2150 & n2818;
  assign n2820 = n2143 & n2819;
  assign n2821 = ~n2131 & n2134;
  assign n2822 = n2146 & ~n2157;
  assign n2823 = ~n2149 & n2822;
  assign n2824 = ~n2153 & n2156;
  assign n2825 = ~n2823 & ~n2824;
  assign n2826 = n2138 & ~n2141;
  assign n2827 = n2825 & ~n2826;
  assign n2828 = n2143 & ~n2827;
  assign n2829 = ~n2821 & ~n2828;
  assign n2830 = ~n2820 & n2829;
  assign n2831 = n2118 & ~n2121;
  assign n2832 = ~n2115 & ~n2831;
  assign n2833 = n2108 & n2832;
  assign n2834 = ~n2830 & n2833;
  assign n2835 = ~n2128 & ~n2834;
  assign n2836 = ~n2126 & n2835;
  assign n2837 = ~n2099 & n2836;
  assign n2838 = \in175  & n1787;
  assign n2839 = \in075  & ~n1787;
  assign n2840 = ~n2838 & ~n2839;
  assign n2841 = \in375  & n1792;
  assign n2842 = \in275  & ~n1792;
  assign n2843 = ~n2841 & ~n2842;
  assign n2844 = n2840 & ~n2843;
  assign n2845 = \in374  & n1792;
  assign n2846 = \in274  & ~n1792;
  assign n2847 = ~n2845 & ~n2846;
  assign n2848 = \in174  & n1787;
  assign n2849 = \in074  & ~n1787;
  assign n2850 = ~n2848 & ~n2849;
  assign n2851 = ~n2847 & n2850;
  assign n2852 = ~n2844 & ~n2851;
  assign n2853 = \in173  & n1787;
  assign n2854 = \in073  & ~n1787;
  assign n2855 = ~n2853 & ~n2854;
  assign n2856 = \in373  & n1792;
  assign n2857 = \in273  & ~n1792;
  assign n2858 = ~n2856 & ~n2857;
  assign n2859 = n2855 & ~n2858;
  assign n2860 = \in372  & n1792;
  assign n2861 = \in272  & ~n1792;
  assign n2862 = ~n2860 & ~n2861;
  assign n2863 = \in172  & n1787;
  assign n2864 = \in072  & ~n1787;
  assign n2865 = ~n2863 & ~n2864;
  assign n2866 = ~n2862 & n2865;
  assign n2867 = ~n2859 & ~n2866;
  assign n2868 = n2852 & n2867;
  assign n2869 = ~n2837 & n2868;
  assign n2870 = ~n2840 & n2843;
  assign n2871 = n2862 & ~n2865;
  assign n2872 = ~n2859 & n2871;
  assign n2873 = ~n2855 & n2858;
  assign n2874 = ~n2872 & ~n2873;
  assign n2875 = n2847 & ~n2850;
  assign n2876 = n2874 & ~n2875;
  assign n2877 = n2852 & ~n2876;
  assign n2878 = ~n2870 & ~n2877;
  assign n2879 = ~n2869 & n2878;
  assign n2880 = n2082 & ~n2085;
  assign n2881 = ~n2079 & ~n2880;
  assign n2882 = n2072 & n2881;
  assign n2883 = ~n2879 & n2882;
  assign n2884 = ~n2092 & ~n2883;
  assign n2885 = ~n2090 & n2884;
  assign n2886 = ~n2063 & n2885;
  assign n2887 = ~n2056 & ~n2886;
  assign n2888 = n2049 & n2887;
  assign n2889 = ~n2034 & n2888;
  assign n2890 = ~n2037 & n2040;
  assign n2891 = n2030 & ~n2056;
  assign n2892 = ~n2033 & n2891;
  assign n2893 = ~n2052 & n2055;
  assign n2894 = ~n2892 & ~n2893;
  assign n2895 = n2044 & ~n2047;
  assign n2896 = n2894 & ~n2895;
  assign n2897 = n2049 & ~n2896;
  assign n2898 = ~n2890 & ~n2897;
  assign n2899 = ~n2889 & n2898;
  assign n2900 = n2017 & ~n2020;
  assign n2901 = ~n2014 & ~n2900;
  assign n2902 = n2007 & n2901;
  assign n2903 = ~n2899 & n2902;
  assign n2904 = ~n2027 & ~n2903;
  assign n2905 = ~n2025 & n2904;
  assign n2906 = ~n1998 & n2905;
  assign n2907 = \in191  & n1787;
  assign n2908 = \in091  & ~n1787;
  assign n2909 = ~n2907 & ~n2908;
  assign n2910 = \in391  & n1792;
  assign n2911 = \in291  & ~n1792;
  assign n2912 = ~n2910 & ~n2911;
  assign n2913 = n2909 & ~n2912;
  assign n2914 = \in390  & n1792;
  assign n2915 = \in290  & ~n1792;
  assign n2916 = ~n2914 & ~n2915;
  assign n2917 = \in190  & n1787;
  assign n2918 = \in090  & ~n1787;
  assign n2919 = ~n2917 & ~n2918;
  assign n2920 = ~n2916 & n2919;
  assign n2921 = ~n2913 & ~n2920;
  assign n2922 = \in189  & n1787;
  assign n2923 = \in089  & ~n1787;
  assign n2924 = ~n2922 & ~n2923;
  assign n2925 = \in389  & n1792;
  assign n2926 = \in289  & ~n1792;
  assign n2927 = ~n2925 & ~n2926;
  assign n2928 = n2924 & ~n2927;
  assign n2929 = \in388  & n1792;
  assign n2930 = \in288  & ~n1792;
  assign n2931 = ~n2929 & ~n2930;
  assign n2932 = \in188  & n1787;
  assign n2933 = \in088  & ~n1787;
  assign n2934 = ~n2932 & ~n2933;
  assign n2935 = ~n2931 & n2934;
  assign n2936 = ~n2928 & ~n2935;
  assign n2937 = n2921 & n2936;
  assign n2938 = ~n2906 & n2937;
  assign n2939 = ~n2909 & n2912;
  assign n2940 = n2931 & ~n2934;
  assign n2941 = ~n2928 & n2940;
  assign n2942 = ~n2924 & n2927;
  assign n2943 = ~n2941 & ~n2942;
  assign n2944 = n2916 & ~n2919;
  assign n2945 = n2943 & ~n2944;
  assign n2946 = n2921 & ~n2945;
  assign n2947 = ~n2939 & ~n2946;
  assign n2948 = ~n2938 & n2947;
  assign n2949 = n1981 & ~n1984;
  assign n2950 = ~n1978 & ~n2949;
  assign n2951 = n1971 & n2950;
  assign n2952 = ~n2948 & n2951;
  assign n2953 = ~n1991 & ~n2952;
  assign n2954 = ~n1989 & n2953;
  assign n2955 = ~n1962 & n2954;
  assign n2956 = ~n1955 & ~n2955;
  assign n2957 = n1948 & n2956;
  assign n2958 = ~n1933 & n2957;
  assign n2959 = ~n1936 & n1939;
  assign n2960 = n1929 & ~n1955;
  assign n2961 = ~n1932 & n2960;
  assign n2962 = ~n1951 & n1954;
  assign n2963 = ~n2961 & ~n2962;
  assign n2964 = n1943 & ~n1946;
  assign n2965 = n2963 & ~n2964;
  assign n2966 = n1948 & ~n2965;
  assign n2967 = ~n2959 & ~n2966;
  assign n2968 = ~n2958 & n2967;
  assign n2969 = n1916 & ~n1919;
  assign n2970 = ~n1913 & ~n2969;
  assign n2971 = n1906 & n2970;
  assign n2972 = ~n2968 & n2971;
  assign n2973 = ~n1926 & ~n2972;
  assign n2974 = ~n1924 & n2973;
  assign n2975 = ~n1897 & n2974;
  assign n2976 = \in1107  & n1787;
  assign n2977 = \in0107  & ~n1787;
  assign n2978 = ~n2976 & ~n2977;
  assign n2979 = \in3107  & n1792;
  assign n2980 = \in2107  & ~n1792;
  assign n2981 = ~n2979 & ~n2980;
  assign n2982 = n2978 & ~n2981;
  assign n2983 = \in3106  & n1792;
  assign n2984 = \in2106  & ~n1792;
  assign n2985 = ~n2983 & ~n2984;
  assign n2986 = \in1106  & n1787;
  assign n2987 = \in0106  & ~n1787;
  assign n2988 = ~n2986 & ~n2987;
  assign n2989 = ~n2985 & n2988;
  assign n2990 = ~n2982 & ~n2989;
  assign n2991 = \in1105  & n1787;
  assign n2992 = \in0105  & ~n1787;
  assign n2993 = ~n2991 & ~n2992;
  assign n2994 = \in3105  & n1792;
  assign n2995 = \in2105  & ~n1792;
  assign n2996 = ~n2994 & ~n2995;
  assign n2997 = n2993 & ~n2996;
  assign n2998 = \in3104  & n1792;
  assign n2999 = \in2104  & ~n1792;
  assign n3000 = ~n2998 & ~n2999;
  assign n3001 = \in1104  & n1787;
  assign n3002 = \in0104  & ~n1787;
  assign n3003 = ~n3001 & ~n3002;
  assign n3004 = ~n3000 & n3003;
  assign n3005 = ~n2997 & ~n3004;
  assign n3006 = n2990 & n3005;
  assign n3007 = ~n2975 & n3006;
  assign n3008 = ~n2978 & n2981;
  assign n3009 = n3000 & ~n3003;
  assign n3010 = ~n2997 & n3009;
  assign n3011 = ~n2993 & n2996;
  assign n3012 = ~n3010 & ~n3011;
  assign n3013 = n2985 & ~n2988;
  assign n3014 = n3012 & ~n3013;
  assign n3015 = n2990 & ~n3014;
  assign n3016 = ~n3008 & ~n3015;
  assign n3017 = ~n3007 & n3016;
  assign n3018 = n1880 & ~n1883;
  assign n3019 = ~n1877 & ~n3018;
  assign n3020 = n1870 & n3019;
  assign n3021 = ~n3017 & n3020;
  assign n3022 = ~n1890 & ~n3021;
  assign n3023 = ~n1888 & n3022;
  assign n3024 = ~n1861 & n3023;
  assign n3025 = ~n1854 & ~n3024;
  assign n3026 = n1847 & n3025;
  assign n3027 = ~n1832 & n3026;
  assign n3028 = ~n1835 & n1838;
  assign n3029 = n1828 & ~n1854;
  assign n3030 = ~n1831 & n3029;
  assign n3031 = ~n1850 & n1853;
  assign n3032 = ~n3030 & ~n3031;
  assign n3033 = n1842 & ~n1845;
  assign n3034 = n3032 & ~n3033;
  assign n3035 = n1847 & ~n3034;
  assign n3036 = ~n3028 & ~n3035;
  assign n3037 = ~n3027 & n3036;
  assign n3038 = n1808 & ~n1818;
  assign n3039 = ~n1815 & ~n3038;
  assign n3040 = n1805 & n3039;
  assign n3041 = ~n3037 & n3040;
  assign n3042 = ~n1825 & ~n3041;
  assign n3043 = ~n1823 & n3042;
  assign n3044 = ~n1796 & n3043;
  assign n3045 = \in1123  & n1787;
  assign n3046 = \in0123  & ~n1787;
  assign n3047 = ~n3045 & ~n3046;
  assign n3048 = \in3123  & n1792;
  assign n3049 = \in2123  & ~n1792;
  assign n3050 = ~n3048 & ~n3049;
  assign n3051 = n3047 & ~n3050;
  assign n3052 = \in3122  & n1792;
  assign n3053 = \in2122  & ~n1792;
  assign n3054 = ~n3052 & ~n3053;
  assign n3055 = \in1122  & n1787;
  assign n3056 = \in0122  & ~n1787;
  assign n3057 = ~n3055 & ~n3056;
  assign n3058 = ~n3054 & n3057;
  assign n3059 = ~n3051 & ~n3058;
  assign n3060 = \in1121  & n1787;
  assign n3061 = \in0121  & ~n1787;
  assign n3062 = ~n3060 & ~n3061;
  assign n3063 = \in3121  & n1792;
  assign n3064 = \in2121  & ~n1792;
  assign n3065 = ~n3063 & ~n3064;
  assign n3066 = n3062 & ~n3065;
  assign n3067 = \in3120  & n1792;
  assign n3068 = \in2120  & ~n1792;
  assign n3069 = ~n3067 & ~n3068;
  assign n3070 = \in1120  & n1787;
  assign n3071 = \in0120  & ~n1787;
  assign n3072 = ~n3070 & ~n3071;
  assign n3073 = ~n3069 & n3072;
  assign n3074 = ~n3066 & ~n3073;
  assign n3075 = n3059 & n3074;
  assign n3076 = ~n3044 & n3075;
  assign n3077 = ~n3047 & n3050;
  assign n3078 = ~n3066 & n3069;
  assign n3079 = ~n3072 & n3078;
  assign n3080 = ~n3062 & n3065;
  assign n3081 = ~n3079 & ~n3080;
  assign n3082 = n3054 & ~n3057;
  assign n3083 = n3081 & ~n3082;
  assign n3084 = n3059 & ~n3083;
  assign n3085 = ~n3077 & ~n3084;
  assign n3086 = ~n3076 & n3085;
  assign n3087 = \in1124  & n1787;
  assign n3088 = \in0124  & ~n1787;
  assign n3089 = ~n3087 & ~n3088;
  assign n3090 = \in3124  & n1792;
  assign n3091 = \in2124  & ~n1792;
  assign n3092 = ~n3090 & ~n3091;
  assign n3093 = n3089 & ~n3092;
  assign n3094 = ~n1213 & n1784;
  assign n3095 = \in1126  & n1787;
  assign n3096 = \in0126  & ~n1787;
  assign n3097 = ~n3095 & ~n3096;
  assign n3098 = \in3126  & n1792;
  assign n3099 = \in2126  & ~n1792;
  assign n3100 = ~n3098 & ~n3099;
  assign n3101 = n3097 & ~n3100;
  assign n3102 = \in1125  & n1787;
  assign n3103 = \in0125  & ~n1787;
  assign n3104 = ~n3102 & ~n3103;
  assign n3105 = \in3125  & n1792;
  assign n3106 = \in2125  & ~n1792;
  assign n3107 = ~n3105 & ~n3106;
  assign n3108 = n3104 & ~n3107;
  assign n3109 = ~n3101 & ~n3108;
  assign n3110 = ~n3094 & n3109;
  assign n3111 = ~n3093 & n3110;
  assign n3112 = ~n3086 & n3111;
  assign n3113 = ~n3089 & n3092;
  assign n3114 = ~n3104 & n3107;
  assign n3115 = ~n3113 & ~n3114;
  assign n3116 = n3109 & ~n3115;
  assign n3117 = ~n3097 & n3100;
  assign n3118 = ~n3116 & ~n3117;
  assign n3119 = ~n3094 & ~n3118;
  assign n3120 = ~n3112 & ~n3119;
  assign \address1  = ~n1785 & n3120;
  assign n3122 = ~n2503 & \address1 ;
  assign n3123 = ~n2500 & ~\address1 ;
  assign \result0  = n3122 | n3123;
  assign n3125 = ~n2497 & \address1 ;
  assign n3126 = ~n2508 & ~\address1 ;
  assign \result1  = n3125 | n3126;
  assign n3128 = ~n2515 & \address1 ;
  assign n3129 = ~n2512 & ~\address1 ;
  assign \result2  = n3128 | n3129;
  assign n3131 = ~n2493 & \address1 ;
  assign n3132 = ~n2490 & ~\address1 ;
  assign \result3  = n3131 | n3132;
  assign n3134 = ~n2484 & \address1 ;
  assign n3135 = ~n2487 & ~\address1 ;
  assign \result4  = n3134 | n3135;
  assign n3137 = ~n2478 & \address1 ;
  assign n3138 = ~n2481 & ~\address1 ;
  assign \result5  = n3137 | n3138;
  assign n3140 = ~n2472 & \address1 ;
  assign n3141 = ~n2475 & ~\address1 ;
  assign \result6  = n3140 | n3141;
  assign n3143 = ~n2468 & \address1 ;
  assign n3144 = ~n2465 & ~\address1 ;
  assign \result7  = n3143 | n3144;
  assign n3146 = ~n2462 & \address1 ;
  assign n3147 = ~n2542 & ~\address1 ;
  assign \result8  = n3146 | n3147;
  assign n3149 = ~n2459 & \address1 ;
  assign n3150 = ~n2549 & ~\address1 ;
  assign \result9  = n3149 | n3150;
  assign n3152 = ~n2455 & \address1 ;
  assign n3153 = ~n2452 & ~\address1 ;
  assign \result10  = n3152 | n3153;
  assign n3155 = ~n2448 & \address1 ;
  assign n3156 = ~n2445 & ~\address1 ;
  assign \result11  = n3155 | n3156;
  assign n3158 = ~n2441 & \address1 ;
  assign n3159 = ~n2438 & ~\address1 ;
  assign \result12  = n3158 | n3159;
  assign n3161 = ~n2434 & \address1 ;
  assign n3162 = ~n2431 & ~\address1 ;
  assign \result13  = n3161 | n3162;
  assign n3164 = ~n2427 & \address1 ;
  assign n3165 = ~n2424 & ~\address1 ;
  assign \result14  = n3164 | n3165;
  assign n3167 = ~n2420 & \address1 ;
  assign n3168 = ~n2417 & ~\address1 ;
  assign \result15  = n3167 | n3168;
  assign n3170 = ~n2414 & \address1 ;
  assign n3171 = ~n2574 & ~\address1 ;
  assign \result16  = n3170 | n3171;
  assign n3173 = ~n2411 & \address1 ;
  assign n3174 = ~n2581 & ~\address1 ;
  assign \result17  = n3173 | n3174;
  assign n3176 = ~n2407 & \address1 ;
  assign n3177 = ~n2404 & ~\address1 ;
  assign \result18  = n3176 | n3177;
  assign n3179 = ~n2400 & \address1 ;
  assign n3180 = ~n2397 & ~\address1 ;
  assign \result19  = n3179 | n3180;
  assign n3182 = ~n2393 & \address1 ;
  assign n3183 = ~n2390 & ~\address1 ;
  assign \result20  = n3182 | n3183;
  assign n3185 = ~n2386 & \address1 ;
  assign n3186 = ~n2383 & ~\address1 ;
  assign \result21  = n3185 | n3186;
  assign n3188 = ~n2379 & \address1 ;
  assign n3189 = ~n2376 & ~\address1 ;
  assign \result22  = n3188 | n3189;
  assign n3191 = ~n2372 & \address1 ;
  assign n3192 = ~n2369 & ~\address1 ;
  assign \result23  = n3191 | n3192;
  assign n3194 = ~n2366 & \address1 ;
  assign n3195 = ~n2606 & ~\address1 ;
  assign \result24  = n3194 | n3195;
  assign n3197 = ~n2363 & \address1 ;
  assign n3198 = ~n2613 & ~\address1 ;
  assign \result25  = n3197 | n3198;
  assign n3200 = ~n2359 & \address1 ;
  assign n3201 = ~n2356 & ~\address1 ;
  assign \result26  = n3200 | n3201;
  assign n3203 = ~n2352 & \address1 ;
  assign n3204 = ~n2349 & ~\address1 ;
  assign \result27  = n3203 | n3204;
  assign n3206 = ~n2345 & \address1 ;
  assign n3207 = ~n2342 & ~\address1 ;
  assign \result28  = n3206 | n3207;
  assign n3209 = ~n2338 & \address1 ;
  assign n3210 = ~n2335 & ~\address1 ;
  assign \result29  = n3209 | n3210;
  assign n3212 = ~n2331 & \address1 ;
  assign n3213 = ~n2328 & ~\address1 ;
  assign \result30  = n3212 | n3213;
  assign n3215 = ~n2324 & \address1 ;
  assign n3216 = ~n2321 & ~\address1 ;
  assign \result31  = n3215 | n3216;
  assign n3218 = ~n2314 & \address1 ;
  assign n3219 = ~n2317 & ~\address1 ;
  assign \result32  = n3218 | n3219;
  assign n3221 = ~n2672 & \address1 ;
  assign n3222 = ~n2669 & ~\address1 ;
  assign \result33  = n3221 | n3222;
  assign n3224 = ~n2683 & \address1 ;
  assign n3225 = ~n2686 & ~\address1 ;
  assign \result34  = n3224 | n3225;
  assign n3227 = ~n2679 & \address1 ;
  assign n3228 = ~n2676 & ~\address1 ;
  assign \result35  = n3227 | n3228;
  assign n3230 = ~n2656 & \address1 ;
  assign n3231 = ~n2653 & ~\address1 ;
  assign \result36  = n3230 | n3231;
  assign n3233 = ~n2663 & \address1 ;
  assign n3234 = ~n2660 & ~\address1 ;
  assign \result37  = n3233 | n3234;
  assign n3236 = ~n2645 & \address1 ;
  assign n3237 = ~n2648 & ~\address1 ;
  assign \result38  = n3236 | n3237;
  assign n3239 = ~n2641 & \address1 ;
  assign n3240 = ~n2638 & ~\address1 ;
  assign \result39  = n3239 | n3240;
  assign n3242 = ~n2295 & \address1 ;
  assign n3243 = ~n2292 & ~\address1 ;
  assign \result40  = n3242 | n3243;
  assign n3245 = ~n2288 & \address1 ;
  assign n3246 = ~n2285 & ~\address1 ;
  assign \result41  = n3245 | n3246;
  assign n3248 = ~n2280 & \address1 ;
  assign n3249 = ~n2277 & ~\address1 ;
  assign \result42  = n3248 | n3249;
  assign n3251 = ~n2272 & \address1 ;
  assign n3252 = ~n2269 & ~\address1 ;
  assign \result43  = n3251 | n3252;
  assign n3254 = ~n2256 & \address1 ;
  assign n3255 = ~n2253 & ~\address1 ;
  assign \result44  = n3254 | n3255;
  assign n3257 = ~n2263 & \address1 ;
  assign n3258 = ~n2260 & ~\address1 ;
  assign \result45  = n3257 | n3258;
  assign n3260 = ~n2245 & \address1 ;
  assign n3261 = ~n2248 & ~\address1 ;
  assign \result46  = n3260 | n3261;
  assign n3263 = ~n2240 & \address1 ;
  assign n3264 = ~n2237 & ~\address1 ;
  assign \result47  = n3263 | n3264;
  assign n3266 = ~n2726 & \address1 ;
  assign n3267 = ~n2729 & ~\address1 ;
  assign \result48  = n3266 | n3267;
  assign n3269 = ~n2767 & \address1 ;
  assign n3270 = ~n2764 & ~\address1 ;
  assign \result49  = n3269 | n3270;
  assign n3272 = ~n2778 & \address1 ;
  assign n3273 = ~n2781 & ~\address1 ;
  assign \result50  = n3272 | n3273;
  assign n3275 = ~n2774 & \address1 ;
  assign n3276 = ~n2771 & ~\address1 ;
  assign \result51  = n3275 | n3276;
  assign n3278 = ~n2755 & \address1 ;
  assign n3279 = ~n2758 & ~\address1 ;
  assign \result52  = n3278 | n3279;
  assign n3281 = ~n2751 & \address1 ;
  assign n3282 = ~n2748 & ~\address1 ;
  assign \result53  = n3281 | n3282;
  assign n3284 = ~n2740 & \address1 ;
  assign n3285 = ~n2743 & ~\address1 ;
  assign \result54  = n3284 | n3285;
  assign n3287 = ~n2736 & \address1 ;
  assign n3288 = ~n2733 & ~\address1 ;
  assign \result55  = n3287 | n3288;
  assign n3290 = ~n2218 & \address1 ;
  assign n3291 = ~n2215 & ~\address1 ;
  assign \result56  = n3290 | n3291;
  assign n3293 = ~n2211 & \address1 ;
  assign n3294 = ~n2208 & ~\address1 ;
  assign \result57  = n3293 | n3294;
  assign n3296 = ~n2203 & \address1 ;
  assign n3297 = ~n2200 & ~\address1 ;
  assign \result58  = n3296 | n3297;
  assign n3299 = ~n2195 & \address1 ;
  assign n3300 = ~n2192 & ~\address1 ;
  assign \result59  = n3299 | n3300;
  assign n3302 = ~n2179 & \address1 ;
  assign n3303 = ~n2176 & ~\address1 ;
  assign \result60  = n3302 | n3303;
  assign n3305 = ~n2186 & \address1 ;
  assign n3306 = ~n2183 & ~\address1 ;
  assign \result61  = n3305 | n3306;
  assign n3308 = ~n2168 & \address1 ;
  assign n3309 = ~n2171 & ~\address1 ;
  assign \result62  = n3308 | n3309;
  assign n3311 = ~n2163 & \address1 ;
  assign n3312 = ~n2160 & ~\address1 ;
  assign \result63  = n3311 | n3312;
  assign n3314 = ~n2146 & \address1 ;
  assign n3315 = ~n2149 & ~\address1 ;
  assign \result64  = n3314 | n3315;
  assign n3317 = ~n2156 & \address1 ;
  assign n3318 = ~n2153 & ~\address1 ;
  assign \result65  = n3317 | n3318;
  assign n3320 = ~n2138 & \address1 ;
  assign n3321 = ~n2141 & ~\address1 ;
  assign \result66  = n3320 | n3321;
  assign n3323 = ~n2134 & \address1 ;
  assign n3324 = ~n2131 & ~\address1 ;
  assign \result67  = n3323 | n3324;
  assign n3326 = ~n2121 & \address1 ;
  assign n3327 = ~n2118 & ~\address1 ;
  assign \result68  = n3326 | n3327;
  assign n3329 = ~n2114 & \address1 ;
  assign n3330 = ~n2111 & ~\address1 ;
  assign \result69  = n3329 | n3330;
  assign n3332 = ~n2103 & \address1 ;
  assign n3333 = ~n2106 & ~\address1 ;
  assign \result70  = n3332 | n3333;
  assign n3335 = ~n2098 & \address1 ;
  assign n3336 = ~n2095 & ~\address1 ;
  assign \result71  = n3335 | n3336;
  assign n3338 = ~n2862 & \address1 ;
  assign n3339 = ~n2865 & ~\address1 ;
  assign \result72  = n3338 | n3339;
  assign n3341 = ~n2858 & \address1 ;
  assign n3342 = ~n2855 & ~\address1 ;
  assign \result73  = n3341 | n3342;
  assign n3344 = ~n2847 & \address1 ;
  assign n3345 = ~n2850 & ~\address1 ;
  assign \result74  = n3344 | n3345;
  assign n3347 = ~n2843 & \address1 ;
  assign n3348 = ~n2840 & ~\address1 ;
  assign \result75  = n3347 | n3348;
  assign n3350 = ~n2085 & \address1 ;
  assign n3351 = ~n2082 & ~\address1 ;
  assign \result76  = n3350 | n3351;
  assign n3353 = ~n2078 & \address1 ;
  assign n3354 = ~n2075 & ~\address1 ;
  assign \result77  = n3353 | n3354;
  assign n3356 = ~n2067 & \address1 ;
  assign n3357 = ~n2070 & ~\address1 ;
  assign \result78  = n3356 | n3357;
  assign n3359 = ~n2062 & \address1 ;
  assign n3360 = ~n2059 & ~\address1 ;
  assign \result79  = n3359 | n3360;
  assign n3362 = ~n2030 & \address1 ;
  assign n3363 = ~n2033 & ~\address1 ;
  assign \result80  = n3362 | n3363;
  assign n3365 = ~n2055 & \address1 ;
  assign n3366 = ~n2052 & ~\address1 ;
  assign \result81  = n3365 | n3366;
  assign n3368 = ~n2044 & \address1 ;
  assign n3369 = ~n2047 & ~\address1 ;
  assign \result82  = n3368 | n3369;
  assign n3371 = ~n2040 & \address1 ;
  assign n3372 = ~n2037 & ~\address1 ;
  assign \result83  = n3371 | n3372;
  assign n3374 = ~n2020 & \address1 ;
  assign n3375 = ~n2017 & ~\address1 ;
  assign \result84  = n3374 | n3375;
  assign n3377 = ~n2013 & \address1 ;
  assign n3378 = ~n2010 & ~\address1 ;
  assign \result85  = n3377 | n3378;
  assign n3380 = ~n2002 & \address1 ;
  assign n3381 = ~n2005 & ~\address1 ;
  assign \result86  = n3380 | n3381;
  assign n3383 = ~n1997 & \address1 ;
  assign n3384 = ~n1994 & ~\address1 ;
  assign \result87  = n3383 | n3384;
  assign n3386 = ~n2931 & \address1 ;
  assign n3387 = ~n2934 & ~\address1 ;
  assign \result88  = n3386 | n3387;
  assign n3389 = ~n2927 & \address1 ;
  assign n3390 = ~n2924 & ~\address1 ;
  assign \result89  = n3389 | n3390;
  assign n3392 = ~n2916 & \address1 ;
  assign n3393 = ~n2919 & ~\address1 ;
  assign \result90  = n3392 | n3393;
  assign n3395 = ~n2912 & \address1 ;
  assign n3396 = ~n2909 & ~\address1 ;
  assign \result91  = n3395 | n3396;
  assign n3398 = ~n1984 & \address1 ;
  assign n3399 = ~n1981 & ~\address1 ;
  assign \result92  = n3398 | n3399;
  assign n3401 = ~n1977 & \address1 ;
  assign n3402 = ~n1974 & ~\address1 ;
  assign \result93  = n3401 | n3402;
  assign n3404 = ~n1966 & \address1 ;
  assign n3405 = ~n1969 & ~\address1 ;
  assign \result94  = n3404 | n3405;
  assign n3407 = ~n1961 & \address1 ;
  assign n3408 = ~n1958 & ~\address1 ;
  assign \result95  = n3407 | n3408;
  assign n3410 = ~n1929 & \address1 ;
  assign n3411 = ~n1932 & ~\address1 ;
  assign \result96  = n3410 | n3411;
  assign n3413 = ~n1954 & \address1 ;
  assign n3414 = ~n1951 & ~\address1 ;
  assign \result97  = n3413 | n3414;
  assign n3416 = ~n1943 & \address1 ;
  assign n3417 = ~n1946 & ~\address1 ;
  assign \result98  = n3416 | n3417;
  assign n3419 = ~n1939 & \address1 ;
  assign n3420 = ~n1936 & ~\address1 ;
  assign \result99  = n3419 | n3420;
  assign n3422 = ~n1919 & \address1 ;
  assign n3423 = ~n1916 & ~\address1 ;
  assign \result100  = n3422 | n3423;
  assign n3425 = ~n1912 & \address1 ;
  assign n3426 = ~n1909 & ~\address1 ;
  assign \result101  = n3425 | n3426;
  assign n3428 = ~n1901 & \address1 ;
  assign n3429 = ~n1904 & ~\address1 ;
  assign \result102  = n3428 | n3429;
  assign n3431 = ~n1896 & \address1 ;
  assign n3432 = ~n1893 & ~\address1 ;
  assign \result103  = n3431 | n3432;
  assign n3434 = ~n3000 & \address1 ;
  assign n3435 = ~n3003 & ~\address1 ;
  assign \result104  = n3434 | n3435;
  assign n3437 = ~n2996 & \address1 ;
  assign n3438 = ~n2993 & ~\address1 ;
  assign \result105  = n3437 | n3438;
  assign n3440 = ~n2985 & \address1 ;
  assign n3441 = ~n2988 & ~\address1 ;
  assign \result106  = n3440 | n3441;
  assign n3443 = ~n2981 & \address1 ;
  assign n3444 = ~n2978 & ~\address1 ;
  assign \result107  = n3443 | n3444;
  assign n3446 = ~n1883 & \address1 ;
  assign n3447 = ~n1880 & ~\address1 ;
  assign \result108  = n3446 | n3447;
  assign n3449 = ~n1876 & \address1 ;
  assign n3450 = ~n1873 & ~\address1 ;
  assign \result109  = n3449 | n3450;
  assign n3452 = ~n1865 & \address1 ;
  assign n3453 = ~n1868 & ~\address1 ;
  assign \result110  = n3452 | n3453;
  assign n3455 = ~n1860 & \address1 ;
  assign n3456 = ~n1857 & ~\address1 ;
  assign \result111  = n3455 | n3456;
  assign n3458 = ~n1828 & \address1 ;
  assign n3459 = ~n1831 & ~\address1 ;
  assign \result112  = n3458 | n3459;
  assign n3461 = ~n1853 & \address1 ;
  assign n3462 = ~n1850 & ~\address1 ;
  assign \result113  = n3461 | n3462;
  assign n3464 = ~n1842 & \address1 ;
  assign n3465 = ~n1845 & ~\address1 ;
  assign \result114  = n3464 | n3465;
  assign n3467 = ~n1838 & \address1 ;
  assign n3468 = ~n1835 & ~\address1 ;
  assign \result115  = n3467 | n3468;
  assign n3470 = ~n1818 & \address1 ;
  assign n3471 = ~n1808 & ~\address1 ;
  assign \result116  = n3470 | n3471;
  assign n3473 = ~n1814 & \address1 ;
  assign n3474 = ~n1811 & ~\address1 ;
  assign \result117  = n3473 | n3474;
  assign n3476 = ~n1800 & \address1 ;
  assign n3477 = ~n1803 & ~\address1 ;
  assign \result118  = n3476 | n3477;
  assign n3479 = ~n1795 & \address1 ;
  assign n3480 = ~n1790 & ~\address1 ;
  assign \result119  = n3479 | n3480;
  assign n3482 = ~n3069 & \address1 ;
  assign n3483 = ~n3072 & ~\address1 ;
  assign \result120  = n3482 | n3483;
  assign n3485 = ~n3065 & \address1 ;
  assign n3486 = ~n3062 & ~\address1 ;
  assign \result121  = n3485 | n3486;
  assign n3488 = ~n3054 & \address1 ;
  assign n3489 = ~n3057 & ~\address1 ;
  assign \result122  = n3488 | n3489;
  assign n3491 = ~n3050 & \address1 ;
  assign n3492 = ~n3047 & ~\address1 ;
  assign \result123  = n3491 | n3492;
  assign n3494 = ~n3092 & \address1 ;
  assign n3495 = ~n3089 & ~\address1 ;
  assign \result124  = n3494 | n3495;
  assign n3497 = ~n3107 & \address1 ;
  assign n3498 = ~n3104 & ~\address1 ;
  assign \result125  = n3497 | n3498;
  assign n3500 = ~n3100 & \address1 ;
  assign n3501 = ~n3097 & ~\address1 ;
  assign \result126  = n3500 | n3501;
  assign n3503 = ~n1213 & n3120;
  assign \result127  = n1784 & ~n3503;
  assign n3505 = n1792 & \address1 ;
  assign n3506 = n1787 & ~\address1 ;
  assign \address0  = n3505 | n3506;
endmodule
