module top (
    \1 , 5, 9, 13, 17, 21, 25, 29, 33, 37, 41, 45, 49, 53, 57, 61, 65, 69,
    73, 77, 81, 85, 89, 93, 97, 101, 105, 109, 113, 117, 121, 125, 129,
    130, 131, 132, 133, 134, 135, 136, 137,
    724, 725, 726, 727, 728, 729, 730, 731, 732, 733, 734, 735, 736, 737,
    738, 739, 740, 741, 742, 743, 744, 745, 746, 747, 748, 749, 750, 751,
    752, 753, 754, 755  );
  input  \1 , 5, 9, 13, 17, 21, 25, 29, 33, 37, 41, 45, 49, 53, 57, 61,
    65, 69, 73, 77, 81, 85, 89, 93, 97, 101, 105, 109, 113, 117, 121, 125,
    129, 130, 131, 132, 133, 134, 135, 136, 137;
  output 724, 725, 726, 727, 728, 729, 730, 731, 732, 733, 734, 735, 736, 737,
    738, 739, 740, 741, 742, 743, 744, 745, 746, 747, 748, 749, 750, 751,
    752, 753, 754, 755;
  wire n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
    n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
    n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113,
    n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
    n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137,
    n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
    n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161,
    n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173,
    n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185,
    n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197,
    n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
    n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
    n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233,
    n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245,
    n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
    n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269,
    n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
    n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293,
    n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305,
    n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317,
    n318, n320, n321, n322, n324, n325, n326, n328, n329, n330, n332, n333,
    n334, n335, n336, n337, n339, n340, n341, n343, n344, n345, n347, n348,
    n349, n351, n352, n353, n354, n355, n356, n357, n359, n360, n361, n363,
    n364, n365, n367, n368, n369, n371, n372, n373, n374, n375, n376, n378,
    n379, n380, n382, n383, n384, n386, n387, n388, n390, n391, n392, n393,
    n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
    n407, n408, n409, n411, n412, n413, n415, n416, n417, n419, n420, n421,
    n422, n423, n425, n426, n427, n429, n430, n431, n433, n434, n435, n437,
    n438, n439, n440, n441, n442, n444, n445, n446, n448, n449, n450, n452,
    n453, n454, n456, n457, n458, n459, n460, n462, n463, n464, n466, n467,
    n468, n470, n471, n472;
  assign n74 = ~\1  & 17;
  assign n75 = \1  & ~17;
  assign n76 = ~n74 & ~n75;
  assign n77 = ~33 & 49;
  assign n78 = 33 & ~49;
  assign n79 = ~n77 & ~n78;
  assign n80 = n76 & ~n79;
  assign n81 = ~n76 & n79;
  assign n82 = ~n80 & ~n81;
  assign n83 = 129 & 137;
  assign n84 = ~65 & 69;
  assign n85 = 65 & ~69;
  assign n86 = ~n84 & ~n85;
  assign n87 = ~73 & 77;
  assign n88 = 73 & ~77;
  assign n89 = ~n87 & ~n88;
  assign n90 = n86 & ~n89;
  assign n91 = ~n86 & n89;
  assign n92 = ~n90 & ~n91;
  assign n93 = ~81 & 85;
  assign n94 = 81 & ~85;
  assign n95 = ~n93 & ~n94;
  assign n96 = ~89 & 93;
  assign n97 = 89 & ~93;
  assign n98 = ~n96 & ~n97;
  assign n99 = n95 & ~n98;
  assign n100 = ~n95 & n98;
  assign n101 = ~n99 & ~n100;
  assign n102 = n92 & ~n101;
  assign n103 = ~n92 & n101;
  assign n104 = ~n102 & ~n103;
  assign n105 = ~n83 & ~n104;
  assign n106 = n83 & n104;
  assign n107 = ~n105 & ~n106;
  assign n108 = n82 & ~n107;
  assign n109 = ~n82 & n107;
  assign n110 = ~n108 & ~n109;
  assign n111 = ~65 & 81;
  assign n112 = 65 & ~81;
  assign n113 = ~n111 & ~n112;
  assign n114 = ~97 & 113;
  assign n115 = 97 & ~113;
  assign n116 = ~n114 & ~n115;
  assign n117 = n113 & ~n116;
  assign n118 = ~n113 & n116;
  assign n119 = ~n117 & ~n118;
  assign n120 = 133 & 137;
  assign n121 = ~\1  & 5;
  assign n122 = \1  & ~5;
  assign n123 = ~n121 & ~n122;
  assign n124 = ~9 & 13;
  assign n125 = 9 & ~13;
  assign n126 = ~n124 & ~n125;
  assign n127 = n123 & ~n126;
  assign n128 = ~n123 & n126;
  assign n129 = ~n127 & ~n128;
  assign n130 = ~17 & 21;
  assign n131 = 17 & ~21;
  assign n132 = ~n130 & ~n131;
  assign n133 = ~25 & 29;
  assign n134 = 25 & ~29;
  assign n135 = ~n133 & ~n134;
  assign n136 = n132 & ~n135;
  assign n137 = ~n132 & n135;
  assign n138 = ~n136 & ~n137;
  assign n139 = n129 & ~n138;
  assign n140 = ~n129 & n138;
  assign n141 = ~n139 & ~n140;
  assign n142 = ~n120 & ~n141;
  assign n143 = n120 & n141;
  assign n144 = ~n142 & ~n143;
  assign n145 = n119 & ~n144;
  assign n146 = ~n119 & n144;
  assign n147 = ~n145 & ~n146;
  assign n148 = ~69 & 85;
  assign n149 = 69 & ~85;
  assign n150 = ~n148 & ~n149;
  assign n151 = ~101 & 117;
  assign n152 = 101 & ~117;
  assign n153 = ~n151 & ~n152;
  assign n154 = n150 & ~n153;
  assign n155 = ~n150 & n153;
  assign n156 = ~n154 & ~n155;
  assign n157 = 134 & 137;
  assign n158 = ~33 & 37;
  assign n159 = 33 & ~37;
  assign n160 = ~n158 & ~n159;
  assign n161 = ~41 & 45;
  assign n162 = 41 & ~45;
  assign n163 = ~n161 & ~n162;
  assign n164 = n160 & ~n163;
  assign n165 = ~n160 & n163;
  assign n166 = ~n164 & ~n165;
  assign n167 = ~49 & 53;
  assign n168 = 49 & ~53;
  assign n169 = ~n167 & ~n168;
  assign n170 = ~57 & 61;
  assign n171 = 57 & ~61;
  assign n172 = ~n170 & ~n171;
  assign n173 = n169 & ~n172;
  assign n174 = ~n169 & n172;
  assign n175 = ~n173 & ~n174;
  assign n176 = n166 & ~n175;
  assign n177 = ~n166 & n175;
  assign n178 = ~n176 & ~n177;
  assign n179 = ~n157 & ~n178;
  assign n180 = n157 & n178;
  assign n181 = ~n179 & ~n180;
  assign n182 = n156 & ~n181;
  assign n183 = ~n156 & n181;
  assign n184 = ~n182 & ~n183;
  assign n185 = ~73 & 89;
  assign n186 = 73 & ~89;
  assign n187 = ~n185 & ~n186;
  assign n188 = ~105 & 121;
  assign n189 = 105 & ~121;
  assign n190 = ~n188 & ~n189;
  assign n191 = n187 & ~n190;
  assign n192 = ~n187 & n190;
  assign n193 = ~n191 & ~n192;
  assign n194 = 135 & 137;
  assign n195 = n129 & ~n166;
  assign n196 = ~n129 & n166;
  assign n197 = ~n195 & ~n196;
  assign n198 = ~n194 & ~n197;
  assign n199 = n194 & n197;
  assign n200 = ~n198 & ~n199;
  assign n201 = n193 & ~n200;
  assign n202 = ~n193 & n200;
  assign n203 = ~n201 & ~n202;
  assign n204 = ~77 & 93;
  assign n205 = 77 & ~93;
  assign n206 = ~n204 & ~n205;
  assign n207 = ~109 & 125;
  assign n208 = 109 & ~125;
  assign n209 = ~n207 & ~n208;
  assign n210 = n206 & ~n209;
  assign n211 = ~n206 & n209;
  assign n212 = ~n210 & ~n211;
  assign n213 = 136 & 137;
  assign n214 = n138 & ~n175;
  assign n215 = ~n138 & n175;
  assign n216 = ~n214 & ~n215;
  assign n217 = ~n213 & ~n216;
  assign n218 = n213 & n216;
  assign n219 = ~n217 & ~n218;
  assign n220 = n212 & ~n219;
  assign n221 = ~n212 & n219;
  assign n222 = ~n220 & ~n221;
  assign n223 = ~5 & 21;
  assign n224 = 5 & ~21;
  assign n225 = ~n223 & ~n224;
  assign n226 = ~37 & 53;
  assign n227 = 37 & ~53;
  assign n228 = ~n226 & ~n227;
  assign n229 = n225 & ~n228;
  assign n230 = ~n225 & n228;
  assign n231 = ~n229 & ~n230;
  assign n232 = 130 & 137;
  assign n233 = ~97 & 101;
  assign n234 = 97 & ~101;
  assign n235 = ~n233 & ~n234;
  assign n236 = ~105 & 109;
  assign n237 = 105 & ~109;
  assign n238 = ~n236 & ~n237;
  assign n239 = n235 & ~n238;
  assign n240 = ~n235 & n238;
  assign n241 = ~n239 & ~n240;
  assign n242 = ~113 & 117;
  assign n243 = 113 & ~117;
  assign n244 = ~n242 & ~n243;
  assign n245 = ~121 & 125;
  assign n246 = 121 & ~125;
  assign n247 = ~n245 & ~n246;
  assign n248 = n244 & ~n247;
  assign n249 = ~n244 & n247;
  assign n250 = ~n248 & ~n249;
  assign n251 = n241 & ~n250;
  assign n252 = ~n241 & n250;
  assign n253 = ~n251 & ~n252;
  assign n254 = ~n232 & ~n253;
  assign n255 = n232 & n253;
  assign n256 = ~n254 & ~n255;
  assign n257 = n231 & ~n256;
  assign n258 = ~n231 & n256;
  assign n259 = ~n257 & ~n258;
  assign n260 = ~9 & 25;
  assign n261 = 9 & ~25;
  assign n262 = ~n260 & ~n261;
  assign n263 = ~41 & 57;
  assign n264 = 41 & ~57;
  assign n265 = ~n263 & ~n264;
  assign n266 = n262 & ~n265;
  assign n267 = ~n262 & n265;
  assign n268 = ~n266 & ~n267;
  assign n269 = 131 & 137;
  assign n270 = n92 & ~n241;
  assign n271 = ~n92 & n241;
  assign n272 = ~n270 & ~n271;
  assign n273 = ~n269 & ~n272;
  assign n274 = n269 & n272;
  assign n275 = ~n273 & ~n274;
  assign n276 = n268 & ~n275;
  assign n277 = ~n268 & n275;
  assign n278 = ~n276 & ~n277;
  assign n279 = ~13 & 29;
  assign n280 = 13 & ~29;
  assign n281 = ~n279 & ~n280;
  assign n282 = ~45 & 61;
  assign n283 = 45 & ~61;
  assign n284 = ~n282 & ~n283;
  assign n285 = n281 & ~n284;
  assign n286 = ~n281 & n284;
  assign n287 = ~n285 & ~n286;
  assign n288 = 132 & 137;
  assign n289 = n101 & ~n250;
  assign n290 = ~n101 & n250;
  assign n291 = ~n289 & ~n290;
  assign n292 = ~n288 & ~n291;
  assign n293 = n288 & n291;
  assign n294 = ~n292 & ~n293;
  assign n295 = n287 & ~n294;
  assign n296 = ~n287 & n294;
  assign n297 = ~n295 & ~n296;
  assign n298 = n110 & n259;
  assign n299 = n278 & n298;
  assign n300 = ~n297 & n299;
  assign n301 = ~n278 & n298;
  assign n302 = n297 & n301;
  assign n303 = n110 & ~n259;
  assign n304 = n278 & n303;
  assign n305 = n297 & n304;
  assign n306 = ~n110 & n259;
  assign n307 = n278 & n306;
  assign n308 = n297 & n307;
  assign n309 = ~n300 & ~n302;
  assign n310 = ~n305 & n309;
  assign n311 = ~n308 & n310;
  assign n312 = ~n147 & n184;
  assign n313 = ~n203 & n312;
  assign n314 = n222 & n313;
  assign n315 = ~n311 & n314;
  assign n316 = ~n110 & n315;
  assign n317 = ~\1  & n316;
  assign n318 = \1  & ~n316;
  assign 724 = n317 | n318;
  assign n320 = ~n259 & n315;
  assign n321 = ~5 & n320;
  assign n322 = 5 & ~n320;
  assign 725 = n321 | n322;
  assign n324 = ~n278 & n315;
  assign n325 = ~9 & n324;
  assign n326 = 9 & ~n324;
  assign 726 = n325 | n326;
  assign n328 = ~n297 & n315;
  assign n329 = ~13 & n328;
  assign n330 = 13 & ~n328;
  assign 727 = n329 | n330;
  assign n332 = n203 & n312;
  assign n333 = ~n222 & n332;
  assign n334 = ~n311 & n333;
  assign n335 = ~n110 & n334;
  assign n336 = ~17 & n335;
  assign n337 = 17 & ~n335;
  assign 728 = n336 | n337;
  assign n339 = ~n259 & n334;
  assign n340 = ~21 & n339;
  assign n341 = 21 & ~n339;
  assign 729 = n340 | n341;
  assign n343 = ~n278 & n334;
  assign n344 = ~25 & n343;
  assign n345 = 25 & ~n343;
  assign 730 = n344 | n345;
  assign n347 = ~n297 & n334;
  assign n348 = ~29 & n347;
  assign n349 = 29 & ~n347;
  assign 731 = n348 | n349;
  assign n351 = n147 & ~n184;
  assign n352 = ~n203 & n351;
  assign n353 = n222 & n352;
  assign n354 = ~n311 & n353;
  assign n355 = ~n110 & n354;
  assign n356 = ~33 & n355;
  assign n357 = 33 & ~n355;
  assign 732 = n356 | n357;
  assign n359 = ~n259 & n354;
  assign n360 = ~37 & n359;
  assign n361 = 37 & ~n359;
  assign 733 = n360 | n361;
  assign n363 = ~n278 & n354;
  assign n364 = ~41 & n363;
  assign n365 = 41 & ~n363;
  assign 734 = n364 | n365;
  assign n367 = ~n297 & n354;
  assign n368 = ~45 & n367;
  assign n369 = 45 & ~n367;
  assign 735 = n368 | n369;
  assign n371 = n203 & n351;
  assign n372 = ~n222 & n371;
  assign n373 = ~n311 & n372;
  assign n374 = ~n110 & n373;
  assign n375 = ~49 & n374;
  assign n376 = 49 & ~n374;
  assign 736 = n375 | n376;
  assign n378 = ~n259 & n373;
  assign n379 = ~53 & n378;
  assign n380 = 53 & ~n378;
  assign 737 = n379 | n380;
  assign n382 = ~n278 & n373;
  assign n383 = ~57 & n382;
  assign n384 = 57 & ~n382;
  assign 738 = n383 | n384;
  assign n386 = ~n297 & n373;
  assign n387 = ~61 & n386;
  assign n388 = 61 & ~n386;
  assign 739 = n387 | n388;
  assign n390 = n147 & n184;
  assign n391 = n203 & n390;
  assign n392 = ~n222 & n391;
  assign n393 = ~n203 & n390;
  assign n394 = n222 & n393;
  assign n395 = n222 & n371;
  assign n396 = n222 & n332;
  assign n397 = ~n392 & ~n394;
  assign n398 = ~n395 & n397;
  assign n399 = ~n396 & n398;
  assign n400 = ~n278 & n306;
  assign n401 = n297 & n400;
  assign n402 = ~n399 & n401;
  assign n403 = ~n147 & n402;
  assign n404 = ~65 & n403;
  assign n405 = 65 & ~n403;
  assign 740 = n404 | n405;
  assign n407 = ~n184 & n402;
  assign n408 = ~69 & n407;
  assign n409 = 69 & ~n407;
  assign 741 = n408 | n409;
  assign n411 = ~n203 & n402;
  assign n412 = ~73 & n411;
  assign n413 = 73 & ~n411;
  assign 742 = n412 | n413;
  assign n415 = ~n222 & n402;
  assign n416 = ~77 & n415;
  assign n417 = 77 & ~n415;
  assign 743 = n416 | n417;
  assign n419 = ~n297 & n307;
  assign n420 = ~n399 & n419;
  assign n421 = ~n147 & n420;
  assign n422 = ~81 & n421;
  assign n423 = 81 & ~n421;
  assign 744 = n422 | n423;
  assign n425 = ~n184 & n420;
  assign n426 = ~85 & n425;
  assign n427 = 85 & ~n425;
  assign 745 = n426 | n427;
  assign n429 = ~n203 & n420;
  assign n430 = ~89 & n429;
  assign n431 = 89 & ~n429;
  assign 746 = n430 | n431;
  assign n433 = ~n222 & n420;
  assign n434 = ~93 & n433;
  assign n435 = 93 & ~n433;
  assign 747 = n434 | n435;
  assign n437 = ~n278 & n303;
  assign n438 = n297 & n437;
  assign n439 = ~n399 & n438;
  assign n440 = ~n147 & n439;
  assign n441 = ~97 & n440;
  assign n442 = 97 & ~n440;
  assign 748 = n441 | n442;
  assign n444 = ~n184 & n439;
  assign n445 = ~101 & n444;
  assign n446 = 101 & ~n444;
  assign 749 = n445 | n446;
  assign n448 = ~n203 & n439;
  assign n449 = ~105 & n448;
  assign n450 = 105 & ~n448;
  assign 750 = n449 | n450;
  assign n452 = ~n222 & n439;
  assign n453 = ~109 & n452;
  assign n454 = 109 & ~n452;
  assign 751 = n453 | n454;
  assign n456 = ~n297 & n304;
  assign n457 = ~n399 & n456;
  assign n458 = ~n147 & n457;
  assign n459 = ~113 & n458;
  assign n460 = 113 & ~n458;
  assign 752 = n459 | n460;
  assign n462 = ~n184 & n457;
  assign n463 = ~117 & n462;
  assign n464 = 117 & ~n462;
  assign 753 = n463 | n464;
  assign n466 = ~n203 & n457;
  assign n467 = ~121 & n466;
  assign n468 = 121 & ~n466;
  assign 754 = n467 | n468;
  assign n470 = ~n222 & n457;
  assign n471 = ~125 & n470;
  assign n472 = 125 & ~n470;
  assign 755 = n471 | n472;
endmodule
